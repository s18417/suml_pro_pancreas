���     �imblearn.pipeline��Pipeline���)��}�(�steps�]�(�maxabsscaler��sklearn.preprocessing._data��MaxAbsScaler���)��}�(�copy���n_features_in_�K�n_samples_seen_�M��max_abs_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����f8�����R�(K�<�NNNJ����J����K t�b�C@     @V@      �?     ��@du��w@i�G5��7@�St$��@ffff&�@    ��@�t�b�scale_�hhK ��h��R�(KK��h �C@     @V@      �?     ��@du��w@i�G5��7@�St$��@ffff&�@    ��@�t�b�_sklearn_version��1.0.1�ub���randomforestclassifier��sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        h,h-ub�n_estimators�Kd�estimator_params�(h;h?h@hAhBhChDhFhEhHt��	bootstrap���	oob_score���n_jobs�NhEK*�verbose�K �
warm_start��hG�balanced��max_samples�Nh;h<h?Nh@KhAKhBG        hC�auto�hDNhFG        hHG        hK�
n_outputs_�K�classes_�hhK ��h��R�(KK��h �C      �?       @      @�t�b�
n_classes_�K�base_estimator_�h9�estimators_�]�(h8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJf��_hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\h�scalar���h�i8�����R�(Kh!NNNJ����J����K t�bC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?K�
node_count�K��nodes�hhK ��h��R�(KK���h�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(h�hlK ��h�hlK��h�hlK��h�h K��h�h K ��h�hlK(��h�h K0��uK8KKt�b�B�(         n                 0]�?*|�m1�?%      �ģR�y}@       e                 �I�f?�^���?�       ���Ǣ2o@       T                 ��\�?����M��?�       Z��F�k@       A                 �k?��	�?w       �e[��f@       >                 `<��?�x�]���?`       ��<-�a@       ;                  �Mm�?���8i�?Y       ӣJ�`@       $                 )DW?]ͤ�?R       �1�|��^@                        �=E?ǂ�Y �?-       �GP�Q@	                        �U��������?%       �G2��L@
                          �P�?���/��?       ���U�5@                        �7�<?�_�A�?
       肵�e`,@                           �?& k�Lj�?       �q��l}@                        T*�
?ʔfm���?       ��Z�N@������������������������       �               ��#���?                         h��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               �k(��"@                        P�$�?��r{��?       e�6� @������������������������       �               ���-��@������������������������       �               ��#���?                        ��"?d6��l�?       ���Aj�A@                        `�]?<&Μ�!�?       D3�\r.@������������������������       �               ���>��@                        � Q	?���/��?       V��7�@������������������������       �               ��/����?                         ��d�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �      �<	       :��,��4@        !                 X?�^�#΀�?       O�{��A%@������������������������       �               �cp>@"       #                 �sM?  k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?%       :                  EHc?�{D���?%       ���YtPK@&       '                 �/��?f�TCA��?"       L����G@������������������������       �               ��#�� @(       3                 �؉�?��-O�?        �����F@)       2                 ���`?"����?        X�[�;@*       -                    �?䱐3+>�?       �'�8�:@+       ,                   Mt? P
�*Q�?       �͉V�M2@������������������������       �               ��#���?������������������������       �               D�JԮD1@.       /                 �ڎ�?�@G���?       hu��@������������������������       �               0����/@0       1                 8לz?z��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               0#0#�?4       5                  �\�?Ԉ�-X�?       q����2@������������������������       �               ��#��@6       9                 �C8�?& k�Lj�?       d*�}#<-@7       8                 $^,W?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@������������������������       �      ��       鰑%@������������������������       �               ���-��@<       =                   ���?ܜ�x�?       d��إV#@������������������������       �               D�JԮD!@������������������������       �      �<       ��#���??       @                 ^�8�?4)�'=P�?        �2"@������������������������       �               ��/����?������������������������       �               0#0# @B       Q                 �[d�?&�R���?       ��y�D@C       F                  �"�?~+"��(�?       �p��6F<@D       E                 ��m\?& k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      �<       ��/���@G       N                 p�7K?��?       |��u�f7@H       I                 �%�q?���cE��?       b�co5@������������������������       �               ��#�� @J       M                  ��?�3���r�?       ��7�nN*@K       L                 pԨ�?�FO���?       �ߌ$@������������������������       �               �k(��"@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       �cp>@O       P                 x5W�?��G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?R       S                  p<��?���Y��?       �m�{��*@������������������������       �               {�5��(@������������������������       �               0#0#�?U       `                 �U:�?Վ�o	�?       -n�JN�B@V       _                  �P�?�*A� f�?       fT�L_4@W       ^                  q�*?rR����?       q\����!@X       Y                    �?�djH�E�?       ^�\m�n@������������������������       �               ��/����?Z       ]                 �R�־L� P?)�?       ����x�@[       \                  @��?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �               �cp>@������������������������       �      ��       \Lg1��&@a       d                  �u��?`�:V��?       �GP�1@b       c                    �?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��	       �P^Cy/@f       m                 0�A�?��Y'Ы�?       �(��*<@g       h                 �=�t?������?       ���y,@������������������������       �               ��#���?i       l                  �~��?�N�+�?       ����*@j       k                    �?|�G���?       ��%�|@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               vb'vb'"@������������������������       �               �C=�C=,@o       �                 ��O�??��3�?�       ̒���k@p                         :��?\����x�?U       O�i��a@q       r                  ��{�?������?       y<���iE@������������������������       �               ��/���@s       x                 �@�?\o��?�?       �>���~C@t       u                 ��^�?z�G���?       '5L�`�'@������������������������       �               ��+��+@v       w                 hJ��?�;�a
=�?       ��l��@������������������������       �               �cp>@������������������������       �               0#0#�?y       z                 `nM�?0�)�n�?       �b�}{.;@������������������������       �               ��+��+4@{       |                 ��޹?d�ih�<�?       ��
@������������������������       �               0#0#@}       ~                 0xP�?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 ��j�?��=�5X�?;       bv���X@�       �                 �&�?�?�0�?9       &�����V@�       �                   �x�?������?       (i�7@�       �                 ���:?hGջ��?       \�W�'3@������������������������       �               �k(��"@�       �                 ����?l�4���?       �tCP��#@������������������������       �               ��/���@�       �                 pč|?z��`p��?       �����@������������������������       �               ��/����?������������������������       �      ��       0#0#@������������������������       �               0����/@�       �                 �ˏ?MR�L�z�?)       ��_���P@�       �                  0Y��?b��$��?       Cb��C@�       �                 PS�~?<�l����?       *s�Q�@@������������������������       �               0#0#@�       �                 8'�?������?       �%Z��;@�       �                 @~��?(r�]i��?       ��U�i�9@�       �                    �?d�r{��?       e�6� @������������������������       �               0����/@�       �                  �?b%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �      ��	       ;l��F:2@������������������������       �               0#0# @�       �                  @���?���!��?       �@��&@�       �                  ��?Ny��]0�?       ���y"@������������������������       �               ��/����?������������������������       �               ��+��+@������������������������       �               ��#���?�       �                 �מp?���?�s�?       �7y}��<@�       �                 ��%�?�y���@�?	       �+�&�G-@�       �                 ��x�?��q�R�?       C}Ԥ@������������������������       �               ��/����?�       �                 P�<�?�J���?       ��*]Y@������������������������       �               0#0# @������������������������       �               ��#�� @������������������������       �      ��       E�JԮD!@�       �                 ��~?      �<	       �C=�C=,@������������������������       �               0#0#�?������������������������       �               ��8��8*@�       �                 0I&�?      �<       �C=�C=@������������������������       �               0#0# @������������������������       �               ��+��+@�       �                  �rm?�<�<.E�?0        2��T@�       �                  c
8? ���'��?       ��1�NA@�       �                 �Z��?���@��?       �<��9@�       �                   �0�?z�G���?       '5L�`�@������������������������       �               �cp>@������������������������       �               H�4H�4@������������������������       �               ��)��)3@�       �                 @�:�?`���?       ��Me�!@�       �                 Ў ]?���WW�?       �j�S@�       �                  ���?�nɵ��?        Cad�J@�       �                  ��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      �<       z�5��@������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �      ��       (S2%S2G@�t�b�values�hhK ��h��R�(KK�KK��h �B�  Gy�5a@鰑Nc@�P��f@Np�}^@�'�xr�V@������C@*���>�]@h
��V@�C=�C=,@�k(���U@]�ڕ��T@��8��8*@-�����K@�+Q��R@#0#0&@-�����K@��z��wR@H�4H�4@�>��nK@Qn��OP@H�4H�4@�GpAF@�e�_��7@        �k(���E@��|��,@        \Lg1��&@鰑%@        <��,��$@��/���@        ��#���?��/���@        ��#���?�cp>@        ��#���?                        �cp>@                ��/����?                ��/����?                ��/����?        �k(��"@                ��#���?���-��@                ���-��@        ��#���?                ���b:@@��/���@        \Lg1��&@��/���@        ���>��@                ��#��@��/���@                ��/����?        ��#��@��/����?                ��/����?        ��#��@                :��,��4@                ��#���?0����/#@                �cp>@        ��#���?��/���@                ��/���@        ��#���?                ;��,��$@�)�B�D@H�4H�4@<��,��$@F�JԮDA@H�4H�4@��#�� @                ��#�� @F�JԮDA@H�4H�4@��#���?�cp>7@H�4H�4@��#���?�cp>7@0#0# @��#���?E�JԮD1@        ��#���?                        D�JԮD1@                �cp>@0#0# @        0����/@                ��/����?0#0# @                0#0# @        ��/����?                        0#0#�?���>��@�cp>'@        ��#��@                z�5��@�cp>'@        z�5��@��/����?                ��/����?        z�5��@                        鰑%@                ���-��@        ��#���?D�JԮD!@                D�JԮD!@        ��#���?                        ��/����?0#0# @        ��/����?                        0#0# @�P^Cy?@D�JԮD!@0#0# @�k(��2@D�JԮD!@0#0#�?��#���?��/���@        ��#���?                        ��/���@        ��,���1@0����/@0#0#�?��,���1@��/���@        ��#�� @                �k(��"@��/���@        �k(��"@��/����?        �k(��"@                        ��/����?                �cp>@                ��/����?0#0#�?                0#0#�?        ��/����?        z�5��(@        0#0#�?{�5��(@                                0#0#�?���b:@@0����/@0#0#�?�P^Cy/@��/���@0#0#�?��#��@��/���@0#0#�?��#��@��/����?0#0#�?        ��/����?        ��#��@        0#0#�?��#�� @        0#0#�?��#�� @                                0#0#�?��#�� @                        �cp>@        \Lg1��&@                ��#��0@��/����?        ��#���?��/����?                ��/����?        ��#���?                �P^Cy/@                ��#���?��/����?k�6k�69@��#���?��/����?#0#0&@��#���?                        ��/����?#0#0&@        ��/����?0#0# @                0#0# @        ��/����?                        vb'vb'"@                �C=�C=,@��#��0@��P@iJ�dJ�a@��b:��*@��|��L@eJ�dJ�Q@        鰑%@0#0#@@        ��/���@                ���-��@0#0#@@        �cp>@H�4H�4@                ��+��+@        �cp>@0#0#�?        �cp>@                        0#0#�?        ��/����?��8��8:@                ��+��+4@        ��/����?H�4H�4@                0#0#@        ��/����?0#0# @        ��/����?                        0#0# @��b:��*@��h
�G@��)��)C@��b:��*@��h
�G@=�C=�C?@�k(��"@鰑%@0#0#@�k(��"@�cp>@0#0#@�k(��"@                        �cp>@0#0#@        ��/���@                ��/����?0#0#@        ��/����?                        0#0#@        0����/@        ��#��@;l��F:B@�;�;;@��#�� @�cp>�9@#0#0&@��#���?��On�8@H�4H�4@                0#0#@��#���?��On�8@0#0# @��#���?��On�8@        ��#���?���-��@                0����/@        ��#���?��/����?                ��/����?        ��#���?                        ;l��F:2@                        0#0# @��#���?��/����?��+��+@        ��/����?��+��+@        ��/����?                        ��+��+@��#���?                ��#�� @鰑%@0#0#0@��#�� @鰑%@0#0# @��#�� @��/����?0#0# @        ��/����?        ��#�� @        0#0# @                0#0# @��#�� @                        E�JԮD!@                        �C=�C=,@                0#0#�?                ��8��8*@                �C=�C=@                0#0# @                ��+��+@z�5��@���-��@gJ�dJ�Q@z�5��@���-��@H�4H�48@        �cp>@#0#06@        �cp>@H�4H�4@        �cp>@                        H�4H�4@                ��)��)3@z�5��@��/���@0#0# @z�5��@��/����?0#0# @z�5��@��/����?0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?z�5��@                                0#0#�?        �cp>@                        (S2%S2G@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�=�KhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKͅ�h��B�,         �                 ���b?f�O?R�?+      \wk]L�}@       �                 0��?�P`��y�?�       +����ku@       ,                 �%{?��n�U�?�       g>Q%�q@       '                 �:W>?^����?M       =��18^@                        �U���\D�R��?B       ��g��*X@                        pe�S?l�R���?       �\���G@                        �-�?l��H��?       ��g���4@������������������������       �               �cp>@	       
                   ��?�Z�	7�?	       ���`�$.@������������������������       �               �cp>@                           �?����?       �Ä�>c(@                        ��?|�6L�n�?       �E#��h @������������������������       �               ��#��@                        ��@?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@                        �Q�?���/��?       V��7�@������������������������       �               ��/����?                         _�
?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?                         ���?��o�G�?       9�� sE9@������������������������       �               ��/����?                         `���?�Wb���?       M�EBCZ7@������������������������       �      ȼ
       z�5��(@                        �N��?�HU����?        ��N��%@                         ���?�_�A�?       肵�e`@������������������������       �               ��/����?������������������������       �               ;��,��@������������������������       �      ��       ��/���@       "                  `�J�?�����?#       ,d�HI@        !                 ;��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?#       $                 p��?�M2�8ӣ?!       i�R�dIH@������������������������       �               ��b:��:@%       &                 pD�\?X ����?       2
C>�5@������������������������       �               ��/����?������������������������       �               <��,��4@(       +                 ����?f��x��?       ̊m68@)       *                  p���?      �<
       鰑5@������������������������       �               ��/���@������������������������       �        	       E�JԮD1@������������������������       �      ȼ       z�5��@-       j                      �n`o4��?n       y>��1�d@.       M                 �[�Z?l�	�<�?B       $�L~VZX@/       :                  �JV�?�z`�m�?       voIi�D@0       7                  ��3�?&���
�?	       䡍�C&@1       6                  �!�?
4=�%�?       �(J��@2       5                 PU1�?Ȕfm���?       ��Z�N@3       4                  kk�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#���?8       9                 PPp�?��ڰ�x�?       �K�f�@������������������������       �               ;��,��@������������������������       �               0#0#�?;       B                  ���?$x����?       ��QR\>@<       =                  P�"�?�֪u�_�?       � Eowj1@������������������������       �               ���-��@>       ?                  `���?������?       +�ǟf%@������������������������       �               0#0#�?@       A                 �m۶?���mf�?       寠�?b#@������������������������       �               0#0# @������������������������       �      ��       ��/���@C       L                  0p��?������?	       Tŵ�)@D       K                  �Mm�?�\`GC��?       � �(&"$@E       J                  �6��?JH����?       ��ϭ
*@F       I                 �_,�?��`i��?       �؛.�@G       H                 �2*�?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?������������������������       �      ȼ       ��/����?������������������������       �               ��#�� @������������������������       �               H�4H�4@������������������������       �      Լ       �cp>@N       a                  I��?�?����?%       ��O���K@O       Z                 �{�?�?�V���?       ���Z~F@P       W                 0�,�?�FO���?       ,��N�>@Q       V                 ��U�?���m�?       ".���<@R       U                 �q�q?X�j���?       ���z"@S       T                 Z��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ��       ���>��@������������������������       �               ������3@X       Y                 �?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?[       \                 �y�?r-�=H�?	       "<��R,@������������������������       �               �k(��"@]       ^                   E(�?���mf�?       毠�?b@������������������������       �               �cp>@_       `                 �Q�?~�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?b       g                 h��? IU����?        ��N��%@c       f                 �j��?�`@s'��?       Ei_y,*@d       e                 �!R�?b%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �               ��/���@h       i                 �=��?      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@k       z                 �F�?R����?,       ��)�FQ@l       s                 ��d�?J���uy�?       v�����6@m       r                 `�*o?��2uj�?	       k溕+@n       q                 �;�?��íxq�?       $2��-�@o       p                 ����?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �      ��       ��/���@������������������������       �               ��/���@t       y                 p?U�?ln����?       ~��Y-"@u       v                  p���?����?       ��X�)B @������������������������       �               ��/����?w       x                 GҎi?l����?       Q	K��@������������������������       �               ��/����?������������������������       �      �<       z�5��@������������������������       �      м       ��/����?{       �                 X�?8s���m�?       k[�ɝ9G@|       �                   ��?��T��u�?       �w8�_@@}       ~                 �V"P?����x�?       �ra6�:@������������������������       �        
       :l��F:2@       �                  ����?�;[��G�?       �O�;�]!@�       �                 艝�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �      �<       ���-��@�       �                  `<��?t@ȱ��?       nm���S@������������������������       �               ��#���?������������������������       �      ��       0����/@�       �                 �j�@?���=�?	       Ԏ{$j+@�       �                 ��E(?�zœ���?       IG���t@������������������������       �               0#0#�?������������������������       �               z�5��@������������������������       �               /����/#@�       �                 �c�?�s�-bS�?#       1�C�K@�       �                 |�L?��OD5�?       �� �D@�       �                 `CN�?�=3��?       �4�zW8@�       �                    �?���­�?	       �##��E0@�       �                  $��?�^h����?       T,��q$@�       �                 p���?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                  9Ρ?��t1u�?       "�te!� @������������������������       �               0#0#�?������������������������       �      ��       ���>��@������������������������       �               H�4H�4@������������������������       �               0#0# @�       �                 �U��?�}h��?       ���r�/@�       �                 �6SZ?��íxq�?	       %2��-�'@�       �                  �d%�?�oH2.w�?       �їD́%@�       �                 ��?�?& k�Lj�?       �q��l}#@������������������������       �               �cp>@�       �                 𡔜?���/��?       V��7�@������������������������       �               ��/����?�       �                 `���?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �               0#0#�?�       �                  c
8?�zœ���?       IG���t@������������������������       �               0#0#�?������������������������       �               z�5��@������������������������       �      ��	       �A�A.@�       �                 Pt%�?P� i���?M       ��R=1`@�       �                  ^�\?fQ ����?       *�_ݗ�#@�       �                  gm?f%@�"�?       ��[�@������������������������       �               ��/����?�       �                 �@�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 ��Խ?�AP�9��?       i��6��@�       �                    �?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0#@�       �                  (��?���Ƚ�?E       ��/���]@�       �                 `�4x?��� ��?0       ux[f��T@�       �                  ;��?��Ñp��?
       ;7��0�%@�       �                 К�?Fy��]0�?       ���y"@�       �                 0��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               0#0#@�       �                 0�2�?���mf�?       毠�?b@������������������������       �               �cp>@�       �                 ���?~�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                    �?H��\ʳ?&       �Q�Fd�Q@������������������������       �               �z��z�B@�       �                 p?�?��Ɵ��?       �(�NA@�       �                  �E�?@�v}�?       ���5>@�       �                   �0�?�n���k�?	       3��&�*@������������������������       �               H�4H�4(@������������������������       �      ȼ       ��/����?������������������������       �               S2%S2%1@�       �                 ���?��G���?       ��%�|@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               �z��z�B@�t�bh�hhK ��h��R�(KK�KK��h �B8  ��b:��c@p�'�x�b@ɔLɔ�d@���khc@�L!��a@8k�6k�G@������a@+����m`@��8��8*@������S@鰑E@        B����R@鰑5@        ��b:��:@/����/3@        �k(��"@�cp>'@                �cp>@        �k(��"@�cp>@                �cp>@        �k(��"@�cp>@        ���>��@��/����?        ��#��@                z�5��@��/����?                ��/����?        z�5��@                ��#�� @��/����?                ��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ��,���1@��/���@                ��/����?        ��,���1@�cp>@        z�5��(@                ;��,��@�cp>@        ;��,��@��/����?                ��/����?        ;��,��@                        ��/���@        6��tSH@��/����?        ��#���?��/����?        ��#���?                        ��/����?        �,����G@��/����?        ��b:��:@                <��,��4@��/����?                ��/����?        <��,��4@                z�5��@鰑5@                鰑5@                ��/���@                E�JԮD1@        z�5��@                ���b:P@���|NV@��8��8*@U^CyeJ@F�JԮDA@��+��+$@<��,��$@h
��6@vb'vb'"@���>��@�cp>@0#0#�?��#�� @�cp>@        ��#���?�cp>@                �cp>@                ��/����?                ��/����?        ��#���?                ��#���?                ;��,��@        0#0#�?;��,��@                                0#0#�?z�5��@1����/3@0#0# @        ��|��,@H�4H�4@        ���-��@                ��/���@H�4H�4@                0#0#�?        ��/���@0#0# @                0#0# @        ��/���@        z�5��@0����/@��+��+@z�5��@��/����?��+��+@z�5��@��/����?0#0# @��#���?��/����?0#0# @��#���?        0#0# @                0#0# @��#���?                        ��/����?        ��#�� @                                H�4H�4@        �cp>@        ���#8E@��On�(@0#0#�?�k(��B@���-��@0#0#�?*�����;@�cp>@        ,�����;@��/����?        ��#�� @��/����?        ��#���?��/����?        ��#���?                        ��/����?        ���>��@                ������3@                        ��/����?                ��/����?                ��/����?        �k(��"@��/���@0#0#�?�k(��"@                        ��/���@0#0#�?        �cp>@                ��/����?0#0#�?                0#0#�?        ��/����?        ;��,��@�cp>@        ��#���?�cp>@        ��#���?��/����?                ��/����?        ��#���?                        ��/���@        ��#��@                ��#���?                z�5��@                ZLg1��&@[�v%jWK@H�4H�4@���>��@��|��,@0#0#�?��#���?�cp>'@0#0#�?��#���?��/���@0#0#�?��#���?        0#0#�?��#���?                                0#0#�?        ��/���@                ��/���@        z�5��@�cp>@        z�5��@��/����?                ��/����?        z�5��@��/����?                ��/����?        z�5��@                        ��/����?        ��#��@&jW�v%D@0#0# @��#���?��/���>@0#0#�?        �cp>�9@0#0#�?        :l��F:2@                ��/���@0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                ���-��@        ��#���?0����/@        ��#���?                        0����/@        z�5��@0����/#@0#0#�?z�5��@        0#0#�?                0#0#�?z�5��@                        /����/#@        z�5��(@D�JԮD!@S2%S2%A@z�5��(@D�JԮD!@��)��)3@���>��@��/����?0#0#0@���>��@��/����?0#0# @���>��@��/����?0#0# @        ��/����?0#0#�?                0#0#�?        ��/����?        ���>��@        0#0#�?                0#0#�?���>��@                                H�4H�4@                0#0# @;��,��@��/���@H�4H�4@��#�� @��/���@0#0# @��#�� @��/���@0#0#�?��#�� @��/���@                �cp>@        ��#�� @��/����?                ��/����?        ��#�� @��/����?        ��#�� @                        ��/����?                        0#0#�?                0#0#�?z�5��@        0#0#�?                0#0#�?z�5��@                                �A�A.@��#���?�cp>'@�s?�s?]@��#���?��/���@��+��+@��#���?��/����?                ��/����?        ��#���?��/����?                ��/����?        ��#���?                        ��/����?��+��+@        ��/����?0#0#�?                0#0#�?        ��/����?                        0#0#@        ��/���@ҷ|˷�[@        ��/���@�z��z�R@        0����/@H�4H�4@        ��/����?��+��+@        ��/����?0#0#�?        ��/����?                        0#0#�?                0#0#@        ��/���@0#0#�?        �cp>@                ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@T2%S2%Q@                �z��z�B@        �cp>@=�C=�C?@        ��/����?�s?�s?=@        ��/����?H�4H�4(@                H�4H�4(@        ��/����?                        S2%S2%1@        ��/����?0#0# @                0#0# @        ��/����?                        �z��z�B@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ\bshFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKՅ�h��B�.         �                 p���?�i��7*�?"      ~' ��l}@       �                 `�2|?F�D�N�?�       �F`M|�t@       D                 ��Ks?�K��{�?�       �ה Er@                        `���?X.����?H       ����8]@                        p|�?�z���`�?       �7���@@                        h7�@?j%@�"�?       Ͱrɱ�=@                        �C[?�HU����?       "��N��5@                           �?d�r{��?       e�6� @	       
                 PO�O?r@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@������������������������       �               ��/����?                         �^��?�f%j��?
       ��ꁞ9,@                        �Q�?�����?	       �Ä�>c(@                        ��aӾ��6L�n�?       �E#��h @                           �?�����?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?������������������������       �               ��#��@                        �@?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      м       ��/����?                        ��Y?      �<       ��/���@������������������������       �               �cp>@������������������������       �               0����/@������������������������       �               ��#��@       +                 �]t?Đ�����?4       �6g�@�T@       $                 �U���L�־+��?!       �I��'3L@       #                 0��j?4=�%�?        �(J��#@                         (�$V?�`@s'��?       Fi_y,*@������������������������       �               ��#���?!       "                 G+�`?      �<       �cp>@������������������������       �               ��/���@������������������������       �               ��/����?������������������������       �      �       z�5��@%       &                 �kd1?�h�xf��?       �)i@G@������������������������       �               Ey�5A@'       *                  `��?xb8�Y�?
       GJͰ(@(       )                 ��c?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               <��,��$@,       5                  ��d�?�<�j���?       vG`���:@-       0                 Е��?�3���r�?	       ��7�nN*@.       /                 `�ռ?      �<       ��#�� @������������������������       �               z�5��@������������������������       �               ;��,��@1       2                 ��;O? k�Lj�?       �q��l}@������������������������       �               �cp>@3       4                 ����?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?6       =                  ��2?D�u7b��?
        ͈��N+@7       :                  �^��?�;[��G�?       �O�;�]!@8       9                 Њ�(?      �<       �cp>@������������������������       �               0����/@������������������������       �               ��/����?;       <                 (�r?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?>       C                 '�Ki?��`i��?       �؛.�@?       B                 `��?D��NV=�?       �t�ܲ@@       A                 0�!�?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               0#0#�?E       \                 Pl֐?����?q       �M(���e@F       [                 P��?@3#܅�?       ���A�@@G       T                 �{`?��|��?       ó�̙4@H       K                  |v?�`@s'��?       Di_y,*+@I       J                 �bu?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?L       O                 pA}?�F���?	       :�.�-'@M       N                 ��?      �<       E�JԮD!@������������������������       �               ��/����?������������������������       �               ���-��@P       S                    �?^%@�"�?       ��[�@Q       R                   �?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      �<       ��/����?U       Z                 P�#�?�)z� ��?       �\�@V       W                  p<��?�d�$���?       �T�f@������������������������       �               ��/����?X       Y                 p�^?      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@������������������������       �      м       ��/����?������������������������       �               ��On�(@]       �                 �^Ҧ?&��&�?Y       ��Mi�a@^       s                 �p�?@�n.��?>       ����X@_       p                  �ni?��H'�@�?       ˿/���H@`       e                 0S�r?�3xO���?       �w�s�iG@a       d                 �$I�?�+�z���?       LGh��
9@b       c                 `bp�?|�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               鰑5@f       i                  �9��?�������?       ݧ�0��5@g       h                  ��~�?d�r{��?       e�6� @������������������������       �               ��#���?������������������������       �               ���-��@j       m                  ���?�.4�v��?	       &�~F�,@k       l                 �1Q?T����?       Q	K��@������������������������       �      �<       z�5��@������������������������       �      ȼ       ��/����?n       o                 �UaG?�w��d��?       �0���s@������������������������       �               H�4H�4@������������������������       �      �<       ��/���@q       r                  ��d�?      �<       H�4H�4@������������������������       �               0#0#�?������������������������       �               0#0# @t       }                 `U�?�
ʭ *�?       Qh�PĶH@u       v                 `q��?.�(��?       ��V-�:@������������������������       �               z�5��(@w       x                 �	�?*�b���?       �GXvƒ,@������������������������       �               ��/����?y       |                 P��?��ڰ�x�?       �K�f�(@z       {                 P���?�J���?       ��*]Y@������������������������       �               ��#�� @������������������������       �               0#0# @������������������������       �      м       ��#�� @~                         �9��?�Z���?       &�K[�6@������������������������       �               0����/@�       �                 ��N�?���cv��?       D��c�1@�       �                  ���?my�|�?
       '�0�-@������������������������       �               ���-��@�       �                 �t��?v��x���?       �!��4 @�       �                 !I�?�_�A�?       肵�e`@�       �                  �G?�?�����?       �O��@������������������������       �      �<       ;��,��@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?������������������������       �               0#0#�?������������������������       �      ȼ       z�5��@�       �                 �v@�?��E@Rm�?       -{�=�E@�       �                 ��?Hy��]0�?       ���y"@������������������������       �               ��/����?������������������������       �               ��+��+@�       �                   �x�?
�*�kH�?       YC�B@�       �                 �t��?h��v���?       7��8@�       �                 P���?$��x1�?       ̓�L2�5@�       �                  �x��?�v���?       ntL�	�1@�       �                 ����?��2uj�?
       l溕+@�       �                 �P��?�+�z���?	       LGh��
)@�       �                 ,���?���mf�?       毠�?b@������������������������       �               0#0#�?������������������������       �      �<       ��/���@������������������������       �               ��/���@������������������������       �      �<       ��#���?�       �                 _%?r�T���?       ��e[�&@�       �                 ,M��?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               0#0#�?�       �                 ��_�?����|e�?       �z �B�@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?������������������������       �               H�4H�4@�       �                    �?      �<       ��On�(@������������������������       �               ��/���@������������������������       �               E�JԮD!@�       �                 �O�?���� ��?       tx[f��D@������������������������       �               �;�;;@�       �                 �/O�?�AP�9��?       h��6��+@�       �                 Ш��?Hy��]0�?       ���y"(@������������������������       �               ��+��+$@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?�       �                 �B�?����n�?R       ��?�Z*a@�       �                 Y�u?&����?5       �Y)��V@������������������������       �               ��/����?�       �                 ��A�?��TZ���?4       c�T13BV@�       �                 0]��?��ݎ3��?1       *{�=�U@�       �                 �qҍ?�u��q�?-       %��<QT@�       �                 �gY�?�$U���?       �}GX�F@�       �                 0�a�?V,�~��?       	s��=;@�       �                 ��N�?��E�B��?       dߞKC.@������������������������       �               ��8��8*@������������������������       �      ȼ       ��/����?�       �                  ;��?�D#���?	       �B�j(@������������������������       �               ��+��+@�       �                 ȮY�?k��9�?       �J���@������������������������       �               H�4H�4@������������������������       �               ��#��@�       �                 pj��?f�*���?
       ���c��1@������������������������       �               ��+��+@�       �                  �G?�?���6�?       0Oi]q)@������������������������       �      ��       E�JԮD!@�       �                 t��I?�J���?       ��*]Y@������������������������       �               ��#�� @������������������������       �               0#0# @������������������������       �               fJ�dJ�A@�       �                 p��?ئ� ��?       rp� k@������������������������       �               ��/���@�       �                 �P��?      �<       0#0# @������������������������       �               0#0#�?������������������������       �               0#0#�?������������������������       �      �       �cp>@�       �                 @�dW?pe�ӔO�?       �R��l/G@�       �                  c
8?����	��?       dR�P�,7@�       �                  P���?�~���9�?       �q�Ί#6@�       �                 �j��?Hy��]0�?       ���y"@������������������������       �               0#0#@�       �                 �qO�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �        	       0#0#0@������������������������       �      �<       ��#���?������������������������       �      ��       %S2%S27@�t�bh�hhK ��h��R�(KK�KK��h �B�  �t�Y,`@Y�ڕ��d@�P�P�e@��>���^@����Xb@2#0#P@��>���^@����-�a@�;�;;@�k(��R@������C@H�4H�4@���>��,@/����/3@        <��,��$@0����/3@        <��,��$@�cp>'@        ��#���?���-��@        ��#���?0����/@        ��#���?                        0����/@                ��/����?        �k(��"@0����/@        �k(��"@�cp>@        ���>��@��/����?        z�5��@��/����?        z�5��@                        ��/����?        ��#��@                ��#�� @��/����?        ��#�� @                        ��/����?                ��/����?                ��/���@                �cp>@                0����/@        ��#��@                Np�}N@%jW�v%4@H�4H�4@~�5��H@���-��@        ��#��@�cp>@        ��#���?�cp>@        ��#���?                        �cp>@                ��/���@                ��/����?        z�5��@                ]Lg1��F@��/����?        Ey�5A@                \Lg1��&@��/����?        ��#���?��/����?                ��/����?        ��#���?                <��,��$@                <��,��$@���-��*@H�4H�4@�k(��"@��/���@        ��#�� @                z�5��@                ;��,��@                ��#���?��/���@                �cp>@        ��#���?��/����?                ��/����?        ��#���?                ��#���?/����/#@H�4H�4@        ��/���@0#0#�?        �cp>@                0����/@                ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?��#���?��/����?0#0# @��#���?��/����?0#0#�?��#���?        0#0#�?                0#0#�?��#���?                        ��/����?                        0#0#�?�,����G@�cp>�Y@H�4H�48@z�5��@���-��:@        z�5��@��|��,@        ��#�� @�cp>'@        ��#���?��/����?                ��/����?        ��#���?                ��#���?鰑%@                E�JԮD!@                ��/����?                ���-��@        ��#���?��/����?        ��#���?��/����?                ��/����?        ��#���?                        ��/����?        ��#��@�cp>@        ��#��@��/����?                ��/����?        ��#��@                ��#���?                z�5��@                        ��/����?                ��On�(@        =��,��D@1����/S@H�4H�48@e:��,&C@��On�H@#0#0&@���>��@F�JԮDA@0#0# @���>��@E�JԮDA@��+��+@        �cp>7@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @        鰑5@        ���>��@�cp>'@H�4H�4@��#���?���-��@        ��#���?                        ���-��@        z�5��@0����/@H�4H�4@z�5��@��/����?        z�5��@                        ��/����?                ��/���@H�4H�4@                H�4H�4@        ��/���@                        H�4H�4@                0#0#�?                0#0# @�P^Cy?@��/���.@H�4H�4@\Lg1��6@��/����?0#0# @z�5��(@                ;��,��$@��/����?0#0# @        ��/����?        <��,��$@        0#0# @��#�� @        0#0# @��#�� @                                0#0# @��#�� @                ��#�� @���-��*@0#0#�?        0����/@        ��#�� @E�JԮD!@0#0#�?;��,��@E�JԮD!@0#0#�?        ���-��@        ;��,��@��/����?0#0#�?;��,��@��/����?        ;��,��@��/����?        ;��,��@                        ��/����?                ��/����?                        0#0#�?z�5��@                z�5��@���-��:@��8��8*@        ��/����?��+��+@        ��/����?                        ��+��+@z�5��@�cp>�9@0#0# @z�5��@���-��*@0#0# @z�5��@���-��*@��+��+@z�5��@��On�(@0#0# @��#���?�cp>'@0#0#�?        �cp>'@0#0#�?        ��/���@0#0#�?                0#0#�?        ��/���@                ��/���@        ��#���?                ��#�� @��/����?0#0#�?��#�� @��/����?        ��#�� @                        ��/����?                        0#0#�?        ��/����?H�4H�4@                H�4H�4@        ��/����?                        H�4H�4@        ��On�(@                ��/���@                E�JԮD!@                ��/���@�z��z�B@                �;�;;@        ��/���@��+��+$@        ��/����?��+��+$@                ��+��+$@        ��/����?                ��/����?        ���>��@&jW�v%4@�����{[@z�5��@1����/3@8��8�cP@        ��/����?        z�5��@E�JԮD1@:��8�cP@z�5��@��|��,@8��8�cP@z�5��@鰑%@N��N��O@z�5��@鰑%@�C=�C=<@��#��@��/����?��-��-5@        ��/����?��8��8*@                ��8��8*@        ��/����?        ��#��@        0#0# @                ��+��+@��#��@        H�4H�4@                H�4H�4@��#��@                ��#�� @D�JԮD!@�C=�C=@                ��+��+@��#�� @E�JԮD!@0#0# @        E�JԮD!@        ��#�� @        0#0# @��#�� @                                0#0# @                fJ�dJ�A@        ��/���@0#0# @        ��/���@                        0#0# @                0#0#�?                0#0#�?        �cp>@        ��#���?��/����?#0#0F@��#���?��/����?��-��-5@        ��/����?��-��-5@        ��/����?��+��+@                0#0#@        ��/����?0#0#�?        ��/����?                        0#0#�?                0#0#0@��#���?                                %S2%S27@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��.hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKυ�h��BH-         �                  b?��B`�;�?)       �7�}@       �                 ����?_&
;8�?�       o��j�v@       t                 ��%~?@�����?�       g��%.r@       K                 P�~�?:Q°�6�?~       � �^{ki@       "                 P�?�*�_�?V       �ͧ��a@                        "?���/��?       ��3�H@                           �?�x�<�?       X&b��q1@                        ��?lb8�Y�?       FJͰ(@	       
                 �K��>�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �               ���>��@                        �v}?�d�$���?       �T�f@������������������������       �               z�5��@                         �JV�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?                        �94W?v+�r7��?       ؖ��<5@@                         �.�?,��c`�?       &��t5)@������������������������       �               ��/���@                        �-�?* k�Lj�?       �q��l}@������������������������       �               �cp>@                        X��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?                        �2�e?$��U>��?       �Y�^�3@������������������������       �               ���>��@                        x��?�L����?       Zk���>)@                           �?f%@�"�?       ��[�@������������������������       �      �<       ��/���@������������������������       �               ��#�� @        !                 �_��?      �<       ���-��@������������������������       �               ��/����?������������������������       �               �cp>@#       ,                 ���5?h�r�-�?7       �FW��V@$       '                  x�>(µ*A
�?
       ��A抌)@%       &                 �K�s?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?(       )                 $��@?" k�Lj�?       �q��l}#@������������������������       �               ��#���?*       +                  ��?�(���?       y��uk!@������������������������       �      �<       ��/���@������������������������       �               ��#���?-       >                 ���@?@o�z�?-       ��L��S@.       =                 �U������f��?!       ���>��M@/       <                 8��?��(���?       �ټ�|=@0       1                 ���T?:d�1s��?       $�!-�=6@������������������������       �               ��/����?2       9                    �?�����?       8�nN�R4@3       8                 Z��?���/��?       V��7�@4       5                 B��g?�d�$���?       �T�f@������������������������       �               ��#�� @6       7                 EĒ?bn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               �cp>@:       ;                 �U�v?lb8�Y�?       FJͰ(@������������������������       �      �<       ZLg1��&@������������������������       �      ȼ       ��/����?������������������������       �               ���>��@������������������������       �               Jp�}>@?       H                 �ڡS?�e�>�?       m�B��3@@       C                 �2OF?���_�?       ���e��#@A       B                 �E��?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?D       E                 ����?�֪u�_�?       ��?�8@������������������������       �               ��/���@F       G                  �"�?z�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?I       J                 P��m?T�j���?       ���z"@������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?L       g                 �m�?�k v|�?(       �J��O@M       Z                 ��Ǆ?LUc��?       ���M�D@N       W                 P�Dv?R^�GH�?       >cmiW6@O       T                 �[q?����?	       ��.�SU-@P       S                 �{q?�}	;	�?       uK�>4%@Q       R                 `�Hj?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               ��/���@U       V                  ���?�����?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?X       Y                  ps�?      �<       ��/���@������������������������       �               ��/����?������������������������       �               ���-��@[       f                 0���?��#���?       �͆�1�2@\       c                  �DN?Jy��]0�?       �N-ۙ2@]       ^                    �?�v�;B��?       ՟���	0@������������������������       �               ��+��+$@_       `                  ��?z��`p��?       �����@������������������������       �               H�4H�4@a       b                 @Ws�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?d       e                 @��?��G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      �<       ��/����?h       o                 Ѐ��?"X���`�?       �� ��4@i       n                  &�Q?޺W�w��?       �'DQm"@j       k                  �jw?u�T���?       ��e[�&@������������������������       �               ��#�� @l       m                �U���?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ;��,��@p       s                 P�s�?t@ȱ��?       nm���S'@q       r                 �ڡS?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      ��       E�JԮD!@u       �                 ���6?(O��r_�?3       B��Ơ�U@v                        @�?خ��p#�?!       R��ҴJO@w       x                 (�_e?|�����?        A{;���N@������������������������       �               ��/����?y       |                     �?|҃l[ �?       Ļ���NN@z       {                  �j?$ k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?}       ~                 `�?.�r?�?       �M�)#�K@������������������������       �               ��b:��J@������������������������       �      �<       ��/����?������������������������       �     ��<       0#0#�?�       �                 ���?_���1�?       d�&v�8@�       �                  
�?¸�qA��?       �����5@�       �                 �D�A?�����?       �O��(@�       �                 ����?f%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �               �k(��"@�       �                 ��k�?�C>�?       �1�m�!@�       �                 pb�?�;�a
=�?       ��l��@�       �                 �M*�?      �<       ��/���@������������������������       �               ��/����?������������������������       �               �cp>@�       �                 �jE?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               ��#�� @�       �                 X��?      �<       ��/���@������������������������       �               ��/����?������������������������       �               �cp>@�       �                  �u��?Lꁘ!O�?/       8*��Q@�       �                 �뜲?�}��3��?&       �h�nwL@�       �                 P���?$�8�4�?       ف��t@@�       �                 0W�?P��~d��?       :E���:@�       �                 `�M�?Z�*z>�?       ����#)@�       �                 ;��?�>s{Ab�?
       `I��n'@�       �                �\Ŗ?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               D�JԮD!@������������������������       �               0#0#�?������������������������       �      �<	       ��|��,@�       �                 PAC�?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0#@�       �                    �?������?       ��8@�       �                 `���?Ǔ�R �?       ��u�(@������������������������       �               �cp>@�       �                  �JV�?���A���?       ��\�F"@������������������������       �      �<       z�5��@�       �                 [x�?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?�       �                 �b\�?Fy��]0�?	       ���y"(@������������������������       �               ��/����?������������������������       �               ��+��+$@�       �                 �+.�?��ih�<�?	       ��
,@�       �                 ��G�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               #0#0&@�       �                 pw\�?�e���?I       ����0�[@�       �                 P�!z?�Qk��?       F�?��4@������������������������       �               0#0# @�       �                  0B�?"@�����?       ]n\�/V)@�       �                 �W�n?��XnP��?       ЭS`oM%@�       �                Z�ϡ?|�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      ȼ       ���-��@������������������������       �               0#0# @�       �                 �K�n?_����?=       ��_�
�V@�       �                  �a�?|��`p��?	       f;3@��1@�       �                 `��?*�Jg@��?       ��G� �%@������������������������       �               ��+��+@������������������������       �               �cp>@������������������������       �               �C=�C=@�       �                 �/O�?�ʊs`�?4       �	S\!R@������������������������       �               �s?�s?=@�       �                 h��?Hc��q��?       �Y�r�E@������������������������       �      ܼ       �;�;;@�       �                 ��? w�;B��?       ՟���	0@������������������������       �               ��/����?�       �                 в��?��(v��?       �A�s(.@������������������������       �               ��+��+$@�       �                  ���?�@����?       ���a�@�       �                  ����?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �      ��       H�4H�4@�t�bh�hhK ��h��R�(KK�KK��h �Bh  )���>bf@�+Q��b@u�qb@)���>bf@����/�`@\��Y��H@���>��e@p%jW�vX@��+��+4@V^CyeZ@h
���S@vb'vb'2@����JW@��h
�G@0#0#�?�#���9@�e�_��7@        �P^Cy/@��/����?        [Lg1��&@��/����?        ��#��@��/����?                ��/����?        ��#��@                ���>��@                ��#��@��/����?        z�5��@                ��#���?��/����?        ��#���?                        ��/����?        <��,��$@h
��6@        ��#���?�cp>'@                ��/���@        ��#���?��/���@                �cp>@        ��#���?��/����?        ��#���?                        ��/����?        �k(��"@鰑%@        ���>��@                ��#�� @鰑%@        ��#�� @��/���@                ��/���@        ��#�� @                        ���-��@                ��/����?                �cp>@        "�}��P@�cp>7@0#0#�?��#��@D�JԮD!@        ��#�� @��/����?        ��#�� @                        ��/����?        ��#�� @��/���@        ��#���?                ��#���?��/���@                ��/���@        ��#���?                $�}��O@��|��,@0#0#�?T^CyeJ@���-��@        ZLg1��6@���-��@        �P^Cy/@���-��@                ��/����?        �P^Cy/@0����/@        ��#��@��/���@        ��#��@��/����?        ��#�� @                ��#�� @��/����?                ��/����?        ��#�� @                        �cp>@        ZLg1��&@��/����?        ZLg1��&@                        ��/����?        ���>��@                Jp�}>@                <��,��$@��/���@0#0#�?��#�� @���-��@0#0#�?��#�� @��/����?        ��#�� @                        ��/����?                0����/@0#0#�?        ��/���@                ��/����?0#0#�?                0#0#�?        ��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        |�5��(@Qn��O@@S2%S2%1@z�5��@h
��6@0#0#0@z�5��@:l��F:2@0#0#�?z�5��@鰑%@0#0#�?        /����/#@0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                ��/���@        z�5��@��/����?        z�5��@                        ��/����?                ��/���@                ��/����?                ���-��@                ��/���@�A�A.@        �cp>@�A�A.@        ��/����?�C=�C=,@                ��+��+$@        ��/����?0#0#@                H�4H�4@        ��/����?0#0#�?                0#0#�?        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?        �k(��"@鰑%@0#0#�?���>��@��/����?0#0#�?��#�� @��/����?0#0#�?��#�� @                        ��/����?0#0#�?        ��/����?                        0#0#�?;��,��@                ��#�� @0����/#@        ��#�� @��/����?        ��#�� @                        ��/����?                E�JԮD!@        "�}��P@;l��F:2@0#0# @�>��nK@���-��@0#0#�?�>��nK@���-��@                ��/����?        �>��nK@�cp>@        ��#���?��/���@                ��/���@        ��#���?                ��b:��J@��/����?        ��b:��J@                        ��/����?                        0#0#�?{�5��(@�cp>'@0#0#�?z�5��(@��/���@0#0#�?<��,��$@��/����?        ��#���?��/����?                ��/����?        ��#���?                �k(��"@                ��#�� @�cp>@0#0#�?        �cp>@0#0#�?        ��/���@                ��/����?                �cp>@                ��/����?0#0#�?                0#0#�?        ��/����?        ��#�� @                        ��/���@                ��/����?                �cp>@        z�5��@����z�A@�s?�s?=@z�5��@�-����@@S2%S2%1@        ���-��:@H�4H�4@        ��On�8@0#0# @        鰑%@0#0# @        鰑%@0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                D�JԮD!@                        0#0#�?        ��|��,@                ��/����?0#0#@        ��/����?                        0#0#@z�5��@���-��@#0#0&@z�5��@0����/@0#0#�?        �cp>@        z�5��@��/����?0#0#�?z�5��@                        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?��+��+$@        ��/����?                        ��+��+$@        ��/����?H�4H�4(@        ��/����?0#0#�?                0#0#�?        ��/����?                        #0#0&@        On��O0@;k�6k�W@        E�JԮD!@H�4H�4(@                0#0# @        E�JԮD!@0#0#@        E�JԮD!@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @        ���-��@                        0#0# @        ��/���@�ڬ�ڬT@        �cp>@H�4H�4(@        �cp>@��+��+@                ��+��+@        �cp>@                        �C=�C=@        ��/����?gJ�dJ�Q@                �s?�s?=@        ��/����?�ڬ�ڬD@                �;�;;@        ��/����?�C=�C=,@        ��/����?                ��/����?�C=�C=,@                ��+��+$@        ��/����?0#0#@        ��/����?0#0#�?                0#0#�?        ��/����?                        H�4H�4@�t�bub�     h,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJj�c;hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK���h��B�&         h                 `<��?Dcx̠O�?      ����.�}@       W                  �/�?�XXK��?�       Y}�]	q@       V                 0!�e?ԍ�VI��?�       +����k@       G                 ���@?�o�A"��?}       ��o|Gj@       2                 ��R�?'T��R��?c       �h	=d@       '                 ~`��9z�J��?F       �⋣˝\@       &                 �I?�ĝ��q�?#       ���^�J@       	                  `s�?�y�8��?       l)�paF@������������������������       �               �cp>@
                           �?���/��?       ��(�D@                        �T?Z��h���?       l��:�=@                         ����?�L����?       Yk���>)@                        �؉�?f%@�"�?       ��[�@������������������������       �               �cp>@                         Pmj�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ��       ���-��@                         p��? r���?       ��|�^1@������������������������       �               ��/����?                         �G?�?��6L�n�?       �E#��h0@                        0� �?k� ѽ?       �����.@                         oEg?T����?       P	K��@������������������������       �               ;��,��@                       �٭�g?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?       %                 ��hn?�4��v�?       �Y-"�'@                          ��g�?x�����?       �4^$4�#@������������������������       �               ��#�� @!       "                 `���>`�r{��?       e�6� @������������������������       �               �cp>@#       $                 h�K?& k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      ��       ��/���@������������������������       �               ��#�� @������������������������       �               ��#�� @(       1                   E(�?|3��F��?#       �V.9�N@)       .                 �6�,? 1_#�?       N!�M<@*       -                    �?�)z� ��?	       `��!5@+       ,                 `?�!?N�ђ���?       �oFݜh%@������������������������       �               ��#�� @������������������������       �      ��       E�JԮD!@������������������������       �               ;��,��$@/       0                 ����>      �<       ���>��@������������������������       �               ��#���?������������������������       �               z�5��@������������������������       �               ��#��@@3       @                 p�Ծ?vT �+��?       ��>Y��G@4       =                 ���x?��3׏O�?       ���W1@@5       6                  ���?�֪u�_�?       ��?�87@������������������������       �               �cp>'@7       8                  ����?�� ��?       qp� k'@������������������������       �               0����/@9       <                    �?�Qk��?       ��Th!�@:       ;                 �X��?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?������������������������       �      �<       ��/����?>       ?                      T���'0�?       �C�� T"@������������������������       �               ���>��@������������������������       �      �<       ��/����?A       F                  �~��?��jN�?	       >@
�.@B       C                 ���?f%@�"�?       ��[�@������������������������       �               ��/����?D       E                 ���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               H�4H�4(@H       K                  �/�?�ݻ�-�?       ��hQ�G@I       J                   +Y�?0���>�?       I�YŦ'5@������������������������       �               $jW�v%4@������������������������       �               0#0#�?L       M                   E(�?x���6��?       �x�I
9@������������������������       �               �cp>@N       Q                    �? s��H��?       �_A�H3@O       P                  ��?�d�$���?       ;��#�.@������������������������       �               z�5��(@������������������������       �      ȼ       �cp>@R       S                  ����?����|e�?       �z �B�@������������������������       �               0#0# @T       U                 0E��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �     ��       �C=�C=,@X       e                 ��<�?�H����?       $
�q.I@Y       d                 P��? �My��?        ��NO,H@Z       c                 p��A?�����?       �O��8@[       \                  ���?L���'0�?       �C�� T2@������������������������       �               ��/����?]       ^                  ��^�?��6L�n�?
       �E#��h0@������������������������       �      �<       ��b:��*@_       `                 x=�?V%@�"�?       ��[�@������������������������       �               ��/����?a       b                 8^7�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               z�5��@������������������������       �               �,����7@f       g                 ��x�?     ��<       0#0# @������������������������       �               0#0#�?������������������������       �               0#0#�?i       �                 �6Sz?�Q����?y       �P"���h@j       �                   p��?*ٓ��?O       �����0`@k       �                 ���?�`��B�?E       ��g�j\@l       �                  �6��?�"��Z��?=       `���Z�X@m       �                 P^��?�:N���?7       �����wV@n       �                 p���?�`֭Q��?2       A�d�@-T@o       �                 ���?��Z�V�?%       �#�7O@p       u                 �>�?ޗ��x$�?       �-�*G@q       t                 �l��?�t����?       b�=�2 @r       s                  �?�����?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?������������������������       �               0#0#@v       y                 �*|}?�`Z#�?       ��8C@w       x                  �jw?b,���O�?       ���/>@������������������������       �               ��#���?������������������������       �               H�4H�4@z       }                    �?��?���?       �c�rA@{       |                 p��?��&���?       ��G2��,@������������������������       �               ���-��*@������������������������       �      �<       ��#���?~                        ��#�?(�ť��?
       7����3@������������������������       �               ��/���@�       �                 �S��?�3`���?       �~�M�(@�       �                 �ss�?�D#���?       ���&P"@�       �                 P�<�?�|2N��?       �3K}@������������������������       �               0#0# @������������������������       �               z�5��@������������������������       �      ��       0#0#@������������������������       �      �<       �cp>@�       �                 @�Ц?�W?Z���?       [�g0@�       �                 �j%?��P����?       <#��,@ @�       �                 ����?�g�vw�?       �Aws}8@�       �                  y��?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               ��#�� @������������������������       �               ��#�� @�       �                 ���?����|e�?       �z �B�@������������������������       �               ��+��+@�       �                 p�)�?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?�       �                 �D��?X,����?       gM��F2@������������������������       �               0#0#�?������������������������       �               D�JԮD1@�       �                 𡔜?R���'0�?       �C�� T"@������������������������       �               ��/����?������������������������       �               ���>��@������������������������       �      ��       D�JԮD!@�       �                  ��?�AP�9��?       i��6��+@������������������������       �               �C=�C=@�       �                 �؉�?�w��d��?       �0���s@������������������������       �               ��/���@������������������������       �      �<       H�4H�4@�       �                 ����?7��b�?
       %�|�1@������������������������       �      ��       ��+��+$@�       �                 ����?X�ih�<�?       ��
@�       �                 �p�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��+��+@�       �                 `�R�?�M��b�?*       7��0��Q@������������������������       �      ȼ       ��-��-E@�       �                  �?`�ih�<�?       ��
<@������������������������       �               ��/����?�       �                 ���?l*�'=P�?       ( AK;@������������������������       �               ��/����?�       �                  ��d�?�n���k�?       3��&�:@�       �                  P�"�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               %S2%S27@�t�bh�hhK ��h��R�(KK�KK��h �B�  cCy��d@Q��+c@�LɔL	c@�#���b@h
��V@vb'vb'B@�#���Y@鰑U@S2%S2%A@�#���Y@鰑U@��+��+4@_Lg1��V@Z�v%jWK@0#0#0@>��,��T@�]�ڕ�?@        Lp�}>@�cp>7@        �k(���5@�cp>7@                �cp>@        �k(���5@&jW�v%4@        ��#��0@���-��*@        ��#�� @鰑%@        ��#�� @��/���@                �cp>@        ��#�� @��/����?                ��/����?        ��#�� @                        ���-��@        ���>��,@�cp>@                ��/����?        ���>��,@��/����?        ���>��,@��/����?        z�5��@��/����?        ;��,��@                ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                        ��/����?        ;��,��@���-��@        z�5��@���-��@        ��#�� @                ��#���?���-��@                �cp>@        ��#���?��/���@        ��#���?                        ��/���@        ��#�� @                ��#�� @                T^CyeJ@E�JԮD!@        ������3@E�JԮD!@        |�5��(@E�JԮD!@        ��#�� @E�JԮD!@        ��#�� @                        E�JԮD!@        ;��,��$@                ���>��@                ��#���?                z�5��@                ��#��@@                ��#�� @�cp>7@0#0#0@���>��@鰑5@0#0#@        0����/3@0#0#@        �cp>'@                ��/���@0#0#@        0����/@                �cp>@0#0#@        ��/����?0#0#@                0#0#@        ��/����?                ��/����?        ���>��@��/����?        ���>��@                        ��/����?        ��#���?��/����?H�4H�4(@��#���?��/����?                ��/����?        ��#���?��/����?                ��/����?        ��#���?                                H�4H�4(@z�5��(@�_��e�=@0#0#@        &jW�v%4@0#0#�?        $jW�v%4@                        0#0#�?z�5��(@0����/#@H�4H�4@        �cp>@        z�5��(@��/���@H�4H�4@z�5��(@�cp>@        z�5��(@                        �cp>@                ��/����?H�4H�4@                0#0# @        ��/����?0#0#�?        ��/����?                        0#0#�?                �C=�C=,@�GpAF@��/���@0#0# @�GpAF@��/���@        :��,��4@��/���@        ���>��,@��/���@                ��/����?        ���>��,@��/����?        ��b:��*@                ��#���?��/����?                ��/����?        ��#���?��/����?        ��#���?                        ��/����?        z�5��@                �,����7@                                0#0# @                0#0#�?                0#0#�?������3@��P@��~���\@������3@;��18N@[��Y��H@������3@�_��e�M@B�A�@@������3@�a#6�K@%S2%S27@������3@��h
�G@%S2%S27@{�5��(@�'�xr�F@%S2%S27@z�5��(@�a#6�;@#0#06@��#�� @��On�8@��8��8*@z�5��@��/����?0#0#@z�5��@��/����?        z�5��@                        ��/����?                        0#0#@;��,��@�e�_��7@vb'vb'"@��#���?        H�4H�4@��#���?                                H�4H�4@��#��@�e�_��7@H�4H�4@��#���?���-��*@                ���-��*@        ��#���?                z�5��@鰑%@H�4H�4@        ��/���@        z�5��@�cp>@H�4H�4@z�5��@        H�4H�4@z�5��@        0#0# @                0#0# @z�5��@                                0#0#@        �cp>@        ��#��@�cp>@vb'vb'"@��#��@��/����?H�4H�4@��#�� @��/����?H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@��#�� @                ��#�� @                        ��/����?H�4H�4@                ��+��+@        ��/����?0#0#�?        ��/����?                        0#0#�?        D�JԮD1@0#0#�?                0#0#�?        D�JԮD1@        ���>��@��/����?                ��/����?        ���>��@                        D�JԮD!@                ��/���@��+��+$@                �C=�C=@        ��/���@H�4H�4@        ��/���@                        H�4H�4@        ��/����?0#0#0@                ��+��+$@        ��/����?H�4H�4@        ��/����?0#0#�?        ��/����?                        0#0#�?                ��+��+@        ��/���@B�A�P@                ��-��-E@        ��/���@H�4H�48@        ��/����?                �cp>@H�4H�48@        ��/����?                ��/����?H�4H�48@        ��/����?0#0#�?                0#0#�?        ��/����?                        %S2%S27@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJGԙGhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhMh�hhK ��h��R�(KM��h��B�9         �                 P���?�G$�5�?+      d�2<xo}@                         ��?p_����?      ��Ѓb�z@       ,                 ���p?2��h�?�       9�]VE�j@       )                 ���?�ʚR��?/       Ж�v��Q@                        ����?\e����?-       �~e�vQ@                        \K�?�\�sF��?
       U>��1@                        ڋr
?p�r{��?       e�6� @������������������������       �               ��#���?	       
                 @.��>      �<       ���-��@������������������������       �               ��/����?������������������������       �               �cp>@������������������������       �               �k(��"@       (                 ��R?p,���O�?#       R^CyeJ@                        ���;?(_k���?       $��IE@                        �U������/��?       J9U6�+@                        p�?Ĕfm���?       ��Z�N@������������������������       �      ��       �cp>@������������������������       �               ��#�� @                        ��?�����?       �O��@                        P� ?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#��@       '                 P�5�? }ZWn��?       p����F<@       &                 �r�?����β�?       ��D�=;@       !                 �hp?� ����?       �	��+9@                         ��i?��|��?       ���ĺw@                         ��,?r@ȱ��?       om���S@������������������������       �      �<       ��/���@                        `��D?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#���?"       %                 X��?�O
�*Q�?
       �͉V�M2@#       $                 0��\?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��/���.@������������������������       �      �<       ��#�� @������������������������       �      �<       ��#���?������������������������       �      ȼ       鰑%@*       +                  P���?     ��<       0#0# @������������������������       �               0#0#�?������������������������       �               0#0#�?-       8                  p��?h��@ʅ�?X       ϥ�V�a@.       1                 �&4�?Ј�-X�?       q����2@/       0                 ���f?�����?       ��X�)B @������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?2       7                 0�F�?�^�#΀�?       O�{��A%@3       6                 �\8?fm���?       ��Z�N@4       5                 ��?�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��/����?������������������������       �               ���-��@9       >                 ��$?�pJ����?M       ��$D-�^@:       ;                 �Q�?(k� ѽ?
       �����.@������������������������       �               ���>��@<       =                 @5�>��6L�n�?       �E#��h @������������������������       �               ��/����?������������������������       �      �<       ���>��@?       n                 0?�l6��?C       Tr W�Z@@       W                 �؉�?B�p"�J�?.       ����ES@A       B                 �7?w���%��?       ����4?@������������������������       �               ��/���@C       P                  ���?�\dO��?       ���ur7@D       G                 �\ͥ?�����?       W!��&@E       F                 0��?b,���O�?       ���/>@������������������������       �               ��#���?������������������������       �               H�4H�4@H       I                 Z��e?���q���?       �:-ߩ�@������������������������       �               ��#�� @J       K                    �?����]L�?       N66�ͯ@������������������������       �               ��/����?L       M                 �~�?��q�R�?       C}Ԥ@������������������������       �               ��#���?N       O                 �И�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?Q       R                   ���?��+%�"�?       ��kw��(@������������������������       �               z�5��@S       T                 p�!�?��ڰ�x�?       �K�f�@������������������������       �               z�5��@U       V                  ���?T����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @X       i                  ���?��ϻN�?       ٕ�F@Y       d                  ���?X
TI
u�?       �إV�C@Z       c                    �?��0��5�?       �8���A@[       `                  �P�?(k� ѽ?       �����.@\       ]                 `��u?\����?       P	K��@������������������������       �               ��#��@^       _                 @��y?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @a       b                 p���?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ���>��@������������������������       �        
       ������3@e       h                 ���m?dn����?       � ��w<@f       g                 �Z�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#���?j       m                  塃?��G9�?       ���=A@k       l                 @*��?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               0#0#@o       ~                 ����?>��㲇�?       T;E�?@p       w                  `���?~�����?       2O�6Nv=@q       r                  �x��?p�i�@M�?       ���wzb0@������������������������       �      �<       鰑%@s       v                   �P�?l@ȱ��?       om���S@t       u                 x��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��/���@x       y                  p�:?��?       ��l}�'*@������������������������       �               �cp>@z       }                 �ݓ�?�d�$���?       �T�f$@{       |                 ���?      �<       ��#�� @������������������������       �               z�5��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?������������������������       �               ��#�� @�       �                  �_�?��-O���?�       ��C��j@�       �                   E(�?��
��?�       ��)xE�h@�       �                 P.ģ?(DgM�?&       ���$GO@�       �                 ��1�?$�_s��?       �+^G@�       �                   ҏ�?%��`�?       Ο@��.(@�       �                 ��L?���mf�?       毠�?b@������������������������       �               �cp>@�       �                 ���?~�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      м       ���>��@�       �                 ����?\���j��?       ��ȥA@������������������������       �               �cp>@�       �                 �:��?PxO�gX�?       ����_<@�       �                   .p�?8n֎~�?       �LW��M:@�       �                 �U��>Ɯf�&��?       �UΔK9@�       �                 @�?4=�%�?       �(J��#@�       �                 И"�?Δfm���?       ��Z�N@������������������������       �               ��#���?�       �                 �~��?�`@s'��?       Ei_y,*@������������������������       �               �cp>@�       �                  @��?Ȕfm���?       ��Z�N@�       �                 P�T�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��#�� @�       �                 ���p?����VV�?	       A�R.�.@������������������������       �               ��|��,@������������������������       �               0#0#�?������������������������       �               0#0#�?�       �                  @��?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?�       �                 ��=�?VF�X��?	       .�=k�U0@������������������������       �               ��/����?�       �                 ��s�?�=�Sο?       ����,@������������������������       �               z�5��(@�       �                 (�q�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 `��a?�ʺ �z�?_       -�J|a@�       �                 ��Fq?�ѲUq��?:       -�x1uV@�       �                 �Y`�?	�j#���?"       |�y�VK@�       �                 0��?�([���?       �p���D@�       �                  `s�?d*�'=P�?        �2"@������������������������       �               �C=�C=@�       �                  v��?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                    �?2��N��?       ��5$<D@@�       �                 `���?z� [��?
       ���x��2@�       �                  $��?)���?       T�M��)@�       �                 pW�?\%��̫�?       �@�o#@�       �                 ��F�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               ��/���@������������������������       �      �<       z�5��@������������������������       �               H�4H�4@�       �                 �5�z?�f�T6|�?
       x,*��P+@������������������������       �               ��#���?�       �                 @���?�L����?	       Yk���>)@������������������������       �               0����/#@�       �                 p�,�?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?�       �                  ���?      �<	       ��8��8*@������������������������       �               0#0#�?������������������������       �               H�4H�4(@�       �                 �Nͼ?&����~�?       �rw���@@�       �                 h�B?�E��y�?       O��TI�:@�       �                 p
E�?k�а.�?       ��W�&2@�       �                 ��ߢ?@�h$g�?	       L(#M?�&@������������������������       �               ��#��@�       �                 �Z�?"�b���?       �GXvƒ@�       �                 ��x�?�����?       �O��@�       �                 �am�?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      ��       z�5��@������������������������       �               0#0#�?�       �                  �ݲ?��|��?       ���ĺw@������������������������       �               0����/@������������������������       �               ��#�� @�       �                  `�J�?)���?       y��uk!@�       �                 `�Q�?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               0����/@�       �                 ����?�Qk��?       ��Th!�@������������������������       �               ��/����?�       �                 @� ?�@����?       ���a�@������������������������       �               ��/����?������������������������       �               0#0#@�       �                 0�#�?te�����?%       X��H@�       �                    �?L�b��?#       ���"G@������������������������       �               S2%S2%1@�       �                 p�?�g�\CY�?       B��(=@�       �                 xܜ�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 PbQ�?l*�'=P�?       ) AK;@������������������������       �               vb'vb'"@�       �                 ����?Jy��]0�?       �N-ۙ2@�       �                 �Qz�?����|e�?
       7\@��'@������������������������       �               0#0#@�       �                 p��z?�~�&��?       ?�]��@������������������������       �               ��/����?�       �                  ���?Hy��]0�?       ���y"@������������������������       �               ��+��+@������������������������       �      ȼ       ��/����?������������������������       �               H�4H�4@�       �                 Vո�?D�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 0"�?@w�;B��?       ՟���	0@������������������������       �               ��8��8*@�       �                 �m�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�                       @8��?(�*�^&�?       d$í�D@�       �                 0g��?t��Y���?       ����B@�       �                 @Ȁ�?�Qk��?       ��Th!�@�       �                   E(�?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �               H�4H�4@                       p���?Hf��{�?       ��C&=@                      @1�?��H�&p�?       L^�3��%@                      �O�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0# @������������������������       �               vb'vb'2@������������������������       �      �       �cp>@�t�bh�hhK ��h��R�(KMKK��h �B�  ������c@��~Y/f@Q��N�a@������c@b�ڕ��d@��8��8Z@��G�[@�cp>W@#0#0&@�,����7@�cp>G@0#0# @�,����7@�cp>G@        ;��,��$@���-��@        ��#���?���-��@        ��#���?                        ���-��@                ��/����?                �cp>@        �k(��"@                ��b:��*@������C@        ��b:��*@��|��<@        ���>��@���-��@        ��#�� @�cp>@                �cp>@        ��#�� @                ;��,��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#��@                z�5��@h
��6@        ;��,��@h
��6@        z�5��@h
��6@        ��#�� @0����/@        ��#���?0����/@                ��/���@        ��#���?��/����?                ��/����?        ��#���?                ��#���?                ��#���?D�JԮD1@        ��#���?��/����?        ��#���?                        ��/����?                ��/���.@        ��#�� @                ��#���?                        鰑%@                        0#0# @                0#0#�?                0#0#�?�k(���U@�cp>G@vb'vb'"@���>��@�cp>'@        z�5��@��/����?        z�5��@                        ��/����?        ��#���?0����/#@        ��#���?�cp>@        ��#���?��/����?                ��/����?        ��#���?                        ��/����?                ���-��@        �b:���S@F�JԮDA@vb'vb'"@���>��,@��/����?        ���>��@                ���>��@��/����?                ��/����?        ���>��@                �P^CyMP@�-����@@vb'vb'"@��b:��J@���-��*@vb'vb'"@�P^Cy/@鰑%@��+��+@        ��/���@        �P^Cy/@�cp>@��+��+@��#��@�cp>@0#0#@��#���?        H�4H�4@��#���?                                H�4H�4@z�5��@�cp>@0#0#�?��#�� @                ��#���?�cp>@0#0#�?        ��/����?        ��#���?��/����?0#0#�?��#���?                        ��/����?0#0#�?                0#0#�?        ��/����?        [Lg1��&@        0#0#�?z�5��@                ;��,��@        0#0#�?z�5��@                ��#�� @        0#0#�?                0#0#�?��#�� @                e:��,&C@�cp>@0#0#@�YLg1B@��/����?        Ey�5A@��/����?        ���>��,@��/����?        z�5��@��/����?        ��#��@                ��#�� @��/����?                ��/����?        ��#�� @                ��#�� @                ��#���?                ���>��@                ������3@                ��#�� @��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#���?                ��#�� @��/����?0#0#@��#�� @��/����?                ��/����?        ��#�� @                                0#0#@ZLg1��&@&jW�v%4@        �k(��"@$jW�v%4@        ��#���?��/���.@                鰑%@        ��#���?0����/@        ��#���?��/����?                ��/����?        ��#���?                        ��/���@        ��#�� @0����/@                �cp>@        ��#�� @��/����?        ��#�� @                z�5��@                ;��,��@                        ��/����?        ��#�� @                ����JG@�+Q��R@2��-�rW@����JG@8l��F:R@�6k�6�S@��b:��:@Qn��O@@H�4H�4@��b:��*@�_��e�=@H�4H�4@���>��@��/���@0#0#�?        ��/���@0#0#�?        �cp>@                ��/����?0#0#�?        ��/����?                        0#0#�?���>��@                z�5��@�cp>�9@0#0# @        �cp>@        z�5��@'jW�v%4@0#0# @��#��@&jW�v%4@0#0# @��#��@&jW�v%4@0#0#�?��#��@�cp>@        ��#�� @�cp>@        ��#���?                ��#���?�cp>@                �cp>@        ��#���?�cp>@        ��#���?��/����?        ��#���?                        ��/����?                ��/����?        ��#�� @                        ��|��,@0#0#�?        ��|��,@                        0#0#�?                0#0#�?��#�� @                ��#���?                ��#���?                ��b:��*@�cp>@                ��/����?        ��b:��*@��/����?        z�5��(@                ��#���?��/����?                ��/����?        ��#���?                ������3@'jW�v%D@��)��)S@������3@����z�A@B�A�@@���>��@0����/3@�C=�C=<@���>��@/����/3@�A�A.@        ��/����?0#0# @                �C=�C=@        ��/����?0#0#�?        ��/����?                        0#0#�?���>��@:l��F:2@�C=�C=@��#��@��/���@�C=�C=@��#��@��/���@0#0#�?��#���?��/���@0#0#�?��#���?        0#0#�?��#���?                                0#0#�?        ��/���@        z�5��@                                H�4H�4@z�5��@鰑%@        ��#���?                ��#�� @鰑%@                0����/#@        ��#�� @��/����?        ��#�� @                        ��/����?                        ��8��8*@                0#0#�?                H�4H�4(@{�5��(@On��O0@��+��+@{�5��(@���-��*@0#0#�?\Lg1��&@�cp>@0#0#�?�k(��"@��/����?0#0#�?��#��@                ;��,��@��/����?0#0#�?;��,��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        z�5��@                                0#0#�?��#�� @0����/@                0����/@        ��#�� @                ��#���?��/���@        ��#���?�cp>@        ��#���?                        �cp>@                0����/@                �cp>@0#0#@        ��/����?                ��/����?0#0#@        ��/����?                        0#0#@        0����/@�
��
�E@        ��/���@��-��-E@                S2%S2%1@        ��/���@k�6k�69@        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@H�4H�48@                vb'vb'"@        �cp>@�A�A.@        �cp>@vb'vb'"@                0#0#@        �cp>@��+��+@        ��/����?                ��/����?��+��+@                ��+��+@        ��/����?                        H�4H�4@        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?�C=�C=,@                ��8��8*@        ��/����?0#0#�?                0#0#�?        ��/����?                鰑%@=�C=�C?@        0����/@=�C=�C?@        �cp>@0#0#@        �cp>@0#0#�?                0#0#�?        �cp>@                        H�4H�4@        ��/����?�;�;;@        ��/����?vb'vb'"@        ��/����?0#0#�?                0#0#�?        ��/����?                        0#0# @                vb'vb'2@        �cp>@        �t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��AhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKم�h��Bx/         �                 pY7e?"�O�WA�?0      D���k}@       �                 �D;�?�.�SE�?�       �*uK��u@                          ҏ�?Ӕ���?�       �XT>�qu@                        �a{?4�|�5�?!       ����^E@                        �t?b%@�"�?       ̰rɱ�-@                          ��?R�ђ���?       �oFݜh%@       
                 �-�? ܜ�x�?
       c��إV#@       	                 ��w�?$ k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?������������������������       �               0����/@������������������������       �      ܼ       ��#���?                         `Lվ����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@                        �T��?  �'1��?       %�B��;@������������������������       �               ���-��*@                        �5R�?t���A�?       0gX\-@������������������������       �               ��#���?                        0�~�?e��}�?
       ��Se+@                        p���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               �cp>'@       �                 ��C?�,M�N]�?�       ���	�r@       �                 p��?�$��n�?�       L�v�zn@       $                 ���U?�*v�o[�?�       C]yQ�9m@       !                 ����?�(�����?	       ��0��0@                         �y����d�$���?       �T�f@                         �P��?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               ��#�� @"       #                    �?      �<       �cp>'@������������������������       �               �cp>@������������������������       �               �cp>@%       :                   Mt?��<7�?�       �~h��%k@&       /                 �U���� �?��?*       q��؆�R@'       ,                 ��V?Fͻ�&��?       {���g�1@(       +                 G+�`?�ۜ�x�?       d��إV#@)       *                 �8`?p�r{��?       e�6� @������������������������       �               ��#���?������������������������       �      ��       ���-��@������������������������       �               ��/����?-       .                 ��=�?����?       ��X�)B @������������������������       �               z�5��@������������������������       �      ȼ       ��/����?0       3                  Ӳ?��G�n�?       ����<L@1       2                 `xNv?����?       ��X�)B0@������������������������       �      ��       {�5��(@������������������������       �      �<       ��/���@4       5                 �$I�?���1�B�?       [����D@������������������������       �               ��/����?6       7                 ��py?P�$3�i�?       ��7���C@������������������������       �               ��,���A@8       9                  �x��?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@;       N                 @ߎ|?�i��?[       �,?/�a@<       M                 0C�?Ӳ(�b��?       .�}Cb;@=       B                    �?�����?       8�nN�R4@>       ?                 `s5�?��t� �?       ����x&@������������������������       �               ;��,��@@       A                 P��?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#��@C       L                 ��V�?Zn����?       ~��Y-"@D       K                 x�9r?�)z� ��?       �\�@E       J                 ����?
4=�%�?       �(J��@F       G                 x��?Δfm���?       ��Z�N@������������������������       �               ��#���?H       I                 g�a?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �               ��#�� @������������������������       �               �C=�C=@O       `                 �h�?vx����?J       ��D-��\@P       U                  ���?�zH3�?       +��Z�9@Q       T                 ��
�?���mf�?       �qB_-@R       S                  �9��?�+�z���?       LGh��
)@������������������������       �               0#0#�?������������������������       �               �cp>'@������������������������       �               0#0# @V       ]                  ���?,�oI���?       ~�V&@W       X                  �Ԧ�?���!��?       �@��&@������������������������       �               ��#���?Y       \                  `���?Ny��]0�?       ���y"@Z       [                   �0�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0#@^       _                 @�ո?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?a       f                  �\�??Mk۪�?:       ���}V@b       e                   �G�?X�j���?       ���z"@c       d                  �/�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               z�5��@g       �                 `�E�?�Ρ����?5       4���i.T@h                          ���?���2��?(       �e9+EBM@i       j                 p'v�?>�]��?       �V�-�@@������������������������       �               ��#�� @k       |                 ���@?;�'��?       F��V�S?@l       {                 ��B�?Ȕfm���?       �2Wd;@m       t                  @V��?j%@�"�?       \��/�4@n       s                   .p�?�_�A�?       肵�e`@o       p                   ��?f%@�"�?       ��[�@������������������������       �               ��/����?q       r                 �=��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#��@u       v                  �~��?�`@s'��?	       Ei_y,*+@������������������������       �               0����/#@w       x                 ��d?���/��?       V��7�@������������������������       �               ��/����?y       z                 �̄�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               ���-��@}       ~                 4�^�?z�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @�       �                  ����?�Z�	7�?       .��9@�       �                 Aј?�FO���?       �ߌ$@�       �                 �N��?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               ���>��@�       �                 P��?4=�%�?       t=�x�-@�       �                 h���?�Z�	7�?	       i~���$@�       �                 ��N�?ʔfm���?       ��Z�N@�       �                  0���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 r��?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?�       �                 �}?�����?       �O��@������������������������       �               ��/����?������������������������       �               ;��,��@������������������������       �      ȼ       0����/@�       �                 PeT�?8���2R�?       _�C�56@������������������������       �               ��+��+@�       �                 ��^�?�S�l�?
       ��8	+*1@�       �                 0Sf�?��íxq�?       $2��-�@�       �                 8�C�?���mf�?       毠�?b@������������������������       �               �cp>@�       �                 X�]�?~�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��#���?�       �                  qm�?D�h$g�?       L(#M?�&@������������������������       �               0#0#�?�       �                 `v"�?�FO���?       �ߌ$@������������������������       �               �k(��"@������������������������       �      ȼ       ��/����?�       �                 �Y�?�?�0�!�?       a`�T�$@������������������������       �               �C=�C=@�       �                  )��?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 @���?D���:�?%       ����EL@�       �                 ���Q?����n8�?$       �:5��3J@�       �                 @Mί?��p�M��?       �$B��A@�       �                 pQ�X?��F���?       ���0�aA@�       �                    �?      �<       E�JԮD1@������������������������       �               E�JԮD!@������������������������       �               E�JԮD!@�       �                    �?r@ȱ��?       ���~1@�       �                 ��_?�O-r��?       �.w��e)@������������������������       �               z�5��@������������������������       �               /����/#@������������������������       �               0����/@������������������������       �      ��       0#0#�?�       �                 �t�?���g��?       �E"zs�0@�       �                ��J;?Iz�9��?
       ��[%@������������������������       �               ��#���?�       �                  `%+�?�5JH���?	       �MOI#@������������������������       �      ��       ��/���@�       �                  �G?�?z�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 �;�?z��`p��?       �����@������������������������       �               0#0#@������������������������       �      �<       ��/����?������������������������       �      �<       ��#��@������������������������       �     ��       H�4H�4@�       �                  ��~�?��Ϙ�?P       R��yfd^@������������������������       �               ��#���?�       �                 �|_�?v=���?O       ,��'"^@�       �                   +Y�?$�0�*�?:       �GU��T@�       �                 � ��?�g���E�?#       �m���I@�       �                 � ̽?H
����?!       ,f�nH@�       �                 @EE�?Xo�k��?        4���G@�       �                 ��{?@�
���?       [��S�B@�       �                  cy?����|e�?       �z �B�@�       �                 P���?X�ih�<�?       ��
@������������������������       �               ��+��+@�       �                 ����?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ȼ       ��/����?������������������������       �      �<       �s?�s?=@�       �                 0���?n��`p��?       f;3@��!@������������������������       �               �cp>@������������������������       �      �<       H�4H�4@������������������������       �      �<       ��/����?�       �                 ��8�?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �               =�C=�C?@������������������������       �               �z��z�B@�t�bh�hhK ��h��R�(KK�KK��h �BX  ��,���a@w�H���e@�dJ�d�c@}�5�wa@�����d@;�;�F@}�5�wa@�����d@������C@���>��@¬��z�A@        ;��,��@/����/#@        ��#�� @D�JԮD!@        ��#���?D�JԮD!@        ��#���?��/���@                ��/���@        ��#���?                        0����/@        ��#���?                z�5��@��/����?                ��/����?        z�5��@                ��#�� @�cp>�9@                ���-��*@        ��#�� @��On�(@        ��#���?                ��#���?��On�(@        ��#���?��/����?                ��/����?        ��#���?                        �cp>'@        ��#��`@��`@������C@�P^Cy_@��]�ڕU@B�A�@@�P^Cy_@�H��tXU@H�4H�48@��#��@��On�(@        ��#��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ��#�� @                        �cp>'@                �cp>@                �cp>@        Np�}^@>l��F:R@H�4H�48@���>��L@On��O0@        ���>��@鰑%@        ��#���?D�JԮD!@        ��#���?���-��@        ��#���?                        ���-��@                ��/����?        z�5��@��/����?        z�5��@                        ��/����?        �}�\I@�cp>@        z�5��(@��/���@        {�5��(@                        ��/���@        e:��,&C@��/����?                ��/����?        e:��,&C@��/����?        ��,���A@                z�5��@��/����?                ��/����?        z�5��@                �P^CyO@P!�ML@H�4H�48@�P^Cy/@0����/@�C=�C=@�P^Cy/@0����/@        �k(��"@��/����?        ;��,��@                ��#��@��/����?                ��/����?        ��#��@                z�5��@�cp>@        ��#��@�cp>@        ��#�� @�cp>@        ��#���?�cp>@        ��#���?                        �cp>@                ��/����?                ��/����?        ��#���?                ��#�� @                ��#�� @                                �C=�C=@����JG@�cp>�I@S2%S2%1@z�5��@��|��,@0#0# @        �cp>'@H�4H�4@        �cp>'@0#0#�?                0#0#�?        �cp>'@                        0#0# @z�5��@�cp>@��+��+@��#���?��/����?��+��+@��#���?                        ��/����?��+��+@        ��/����?0#0#�?                0#0#�?        ��/����?                        0#0#@��#�� @��/����?        ��#�� @                        ��/����?        �k(���E@�+Q��B@vb'vb'"@��#�� @��/����?        ��#�� @��/����?                ��/����?        ��#�� @                z�5��@                ��,���A@<l��F:B@vb'vb'"@~�5��8@�]�ڕ�?@0#0# @�k(��"@h
��6@0#0# @��#�� @                ���>��@h
��6@0#0# @���>��@%jW�v%4@        ���>��@���-��*@        ;��,��@��/����?        ��#���?��/����?                ��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#��@                ��#�� @�cp>'@                0����/#@        ��#�� @��/����?                ��/����?        ��#�� @��/����?                ��/����?        ��#�� @                        ���-��@                ��/����?0#0# @        ��/����?                        0#0# @�P^Cy/@/����/#@        �k(��"@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ���>��@                z�5��@E�JԮD!@        z�5��@��/���@        ��#���?�cp>@        ��#���?��/����?                ��/����?        ��#���?                        ��/����?                ��/����?                ��/����?        ;��,��@��/����?                ��/����?        ;��,��@                        0����/@        <��,��$@0����/@�C=�C=@                ��+��+@;��,��$@0����/@0#0# @��#���?��/���@0#0#�?        ��/���@0#0#�?        �cp>@                ��/����?0#0#�?        ��/����?                        0#0#�?��#���?                �k(��"@��/����?0#0#�?                0#0#�?�k(��"@��/����?        �k(��"@                        ��/����?                ��/����?vb'vb'"@                �C=�C=@        ��/����?0#0# @        ��/����?                        0#0# @��#�� @鰑E@H�4H�4@��#��@鰑E@H�4H�4@z�5��@�]�ڕ�?@0#0#�?z�5��@�]�ڕ�?@                E�JԮD1@                E�JԮD!@                E�JԮD!@        z�5��@��|��,@        z�5��@0����/#@        z�5��@                        /����/#@                0����/@                        0#0#�?��#���?鰑%@��+��+@��#���?D�JԮD!@0#0#�?��#���?                        E�JԮD!@0#0#�?        ��/���@                ��/����?0#0#�?                0#0#�?        ��/����?                ��/����?0#0#@                0#0#@        ��/����?        ��#��@                                H�4H�4@��#���?0����/#@�+��+�[@��#���?                        0����/#@�+��+�[@        0����/#@���~�gR@        /����/#@��-��-E@        ���-��@�ڬ�ڬD@        0����/@�ڬ�ڬD@        ��/����?eJ�dJ�A@        ��/����?H�4H�4@        ��/����?H�4H�4@                ��+��+@        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?                        �s?�s?=@        �cp>@H�4H�4@        �cp>@                        H�4H�4@        ��/����?                �cp>@0#0#�?        �cp>@                        0#0#�?                =�C=�C?@                �z��z�B@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ,�hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK兔h��B2         �                   �0�?��։P�?*      dr� z}@       �                 ��x�?��Sy�<�?�       &���жs@       h                  �/�?f7�c5�?�       KT��.Gr@       %                 ���T?��Ez�?�       ����i@       "                 ��]"?���P#�?1       �fX��S@                         ��d�?�.R����?&       �z���M@                        `%�7?�HU����?!       lgP�.TK@                        @F��)z� ��?       a��!E@	                         =�m?�=����?       6��cxA@
                          �P�?hy8�n�?	       O(�\S'/@                        P���>
��I@�?       �2d�%@������������������������       �               0����/@                         h��?���/��?       Az$S��@������������������������       �               z�5��@                           �?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               0����/@                        X\ ?d�WT�V�?	       D$_]3@                        �^o?      �<       �P^Cy/@������������������������       �               ;��,��@������������������������       �               ;��,��$@������������������������       �      �<       ��/���@                         eE7?d����?       P	K��@������������������������       �               ��/����?������������������������       �               z�5��@                        P>-l?$��c`�?
       $��t5)@������������������������       �      ��	       �cp>'@������������������������       �      �<       ��#���?                        ����?�d�$���?       �T�f@������������������������       �               ��/����?        !                 �$?      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@#       $                ��x�'?      �<       �k(��2@������������������������       �               ��#���?������������������������       �        
       ��,���1@&       U                 �\�?�bJ`h��?R       �[V!�_@'       6                  �_�?
��8��?:       �Cm��W@(       3                 �4p?*h��g&�?       㚨\�@@)       0                 `�7�? �l���?       ��P:j�3@*       +                 �U�?& k�Lj�?       d*�}#<-@������������������������       �               E�JԮD!@,       -                 �%�C?���/��?       Az$S��@������������������������       �               z�5��@.       /                 @���?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?1       2                  s��?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?4       5                 ���?      �<       ���-��*@������������������������       �               ��/����?������������������������       �               ��On�(@7       P                  �v�?P4�K���?(       '�?��N@8       M                 )��?f%@�"�?        ��[�G@9       D                 ��Yk?4=�%�?       �(J��C@:       ?                  �\�?p@ȱ��?       nm���S7@;       <                 ���N?Bǵ3���?       �q�ͨ�@������������������������       �               z�5��@=       >                    �?      �<       0����/@������������������������       �               �cp>@������������������������       �               ��/����?@       A                 L��R?�Tu��?	       ����.@������������������������       �               �cp>'@B       C                 `9�`?̔fm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@E       L                  �Ԧ�? ����?       ��X�)B0@F       I                 0�?\����?       R	K��,@G       H                 p���>      �<	       �k(��"@������������������������       �               ��#���?������������������������       �               ��#�� @J       K                 4��?֗Z�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@������������������������       �      ȼ       ��/����?N       O                 pl�]?      �<       ��/���@������������������������       �               ��/����?������������������������       �               �cp>@Q       T                 p���?�26�
�?       4��*8E,@R       S                 ��K�?L� P?)�?       ����x�$@������������������������       �               0#0# @������������������������       �               ��#�� @������������������������       �      ȼ       ��/���@V       g                 ��?�I=8�?       ����<R@@W       f                 p���?p2'��?       �����8@X       a                 �O�?�{�M���?       ��?8�4@Y       Z                 h�B?*^�yU�?	       ��7�1�#@������������������������       �               0#0#@[       \                 p���?x�G���?       '5L�`�@������������������������       �               ��/����?]       ^                 <�Q?����|e�?       �z �B�@������������������������       �               0#0# @_       `                 [�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?b       e                 `��?�}	;	�?       vK�>4%@c       d                 ʎ ]?���mf�?       毠�?b@������������������������       �      �<       ��/���@������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �               0#0#@������������������������       �               0#0# @i       ~                 ��?�c�ms��?0       �����U@j       u                 pW��?�q��j��?        �r`�k�N@k       t                 �U:�?�v^�n�?       ��m�G@l       m                 �5%?�o����?       ���5u:@������������������������       �               ��#��0@n       q                 �n�?4=�%�?       �(J��#@o       p                 ��q?�`@s'��?       Ei_y,*@������������������������       �               ��#���?������������������������       �               �cp>@r       s                    �?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �        	       <��,��4@v       }                  (��?��z�?	       ������,@w       |                 P��?��oR��?       l�Q6�(@x       y                 ���?|���X��?       &��֞&@������������������������       �               �k(��"@z       {                 �jE?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �               0#0# @       �                   E(�?@���v�?       �V��{9@������������������������       �               D�JԮD!@�       �                    �?�K����?       C1��0@�       �                 @�>�?~�G���?       (5L�`�'@�       �                  ��?<�a
=�?       ��l��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �               ��+��+@������������������������       �               ��+��+@�       �                   ���?6��5r�?       ��#�%�6@������������������������       �               �C=�C=@�       �                  �\�?��B��?       sy(��/@������������������������       �               ��/����?�       �                 �y�?���b�?
       �{u;y�-@������������������������       �               ��#���?�       �                  �/�?�AP�9��?	       h��6��+@������������������������       �               ��/����?�       �                   s��?Hy��]0�?       ���y"(@�       �                 ����?lutee�?       Q9��@�       �                 0翇?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0# @������������������������       �      ��       �C=�C=@�       �                 �U,�?����Y�?i       �ʝ���c@�       �                 Џ�b?�!�|��?"       #�h�ГF@�       �                 ��΢?��t�%��?       �u�XD@�       �                  �Mm�?fn����?       րh��K>@�       �                 `8X?�����?       8�nN�R4@������������������������       �               ��/����?�       �                 �R3|?b�WT�V�?       D$_]3@�       �                 ��'�?xb8�Y�?	       FJͰ(@������������������������       �               ;��,��$@�       �                 �/��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 �3?�)z� ��?       �\�@������������������������       �               �cp>@������������������������       �               ��#��@�       �                  �?���/��?       5��o��#@�       �                 �~�?$ k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      ��       ��/���@�       �                 0I��?�d�$���?       �T�f@�       �                  b��>      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@������������������������       �      ȼ       ��/����?�       �                 p�?l?Z@ �F��?       uռ7�#@�       �                 ����?lutee�?       Q9��@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?�       �                    �?* k�Lj�?       �q��l}@�       �                 0�Q�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                  ,�f?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?�       �                 �Ҵn?      �<       ��+��+@������������������������       �               0#0#�?������������������������       �               0#0#@�       �                  �fq?���.1��?G       �V�[@�       �                 �I��?���!��?'       ��{�1XL@�       �                   Y��?;.as���?       =�J�2�C@�       �                 0/|�?�Y�Z�?       X�S��u;@�       �                  `���?� ����?       J���/@�       �                 Yש�?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?�       �                 �u��?�ڇ���?
       4Y����'@������������������������       �               �cp>@�       �                 �8�?�4^��?       s_w$/"@�       �                 �۶�?��q�R�?       B}Ԥ@�       �                 �25�?x�G���?       ��%�|@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �               H�4H�4@�       �                ��2yt?�>s{Ab�?       aI��n'@������������������������       �               0#0#�?������������������������       �               鰑%@�       �                 H<��?��]ۀ��?	       F���O(@������������������������       �               ��#���?�       �                 �]��?���3�?       &��X&@�       �                  ��?޾�R���?       :�S) $@�       �                 (��?X*�'=P�?        �2"@������������������������       �               ��+��+@�       �                 0�H�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �      �<       ��#���?������������������������       �      ȼ       ��/����?�       �                 �둗?(,N=� �?       ��a��+1@������������������������       �        	       �C=�C=,@�       �                 ����?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?�       �                  N��?p�)�n�?        �b�}{.K@������������������������       �               ��-��-E@�       �                 ����?Py��]0�?       ���y"(@������������������������       �               ��/����?������������������������       �               ��+��+$@�t�b�d     h�hhK ��h��R�(KK�KK��h �Bx  �����c@�)�B�d@�4H�4�b@�t�Y,`@��`@�[��[�L@���b:`@k>�c�^@��+��+D@f:��,&S@(�B��Y@��8��8:@6��tSH@�_��e�=@        Lp�}>@�_��e�=@        
�#���9@��|��<@        |�5��8@D�JԮD1@        �k(��2@On��O0@        z�5��@��On�(@        z�5��@��/���@                0����/@        z�5��@�cp>@        z�5��@                        �cp>@                ��/����?                ��/����?                0����/@        �P^Cy/@��/���@        �P^Cy/@                ;��,��@                ;��,��$@                        ��/���@        z�5��@��/����?                ��/����?        z�5��@                ��#���?�cp>'@                �cp>'@        ��#���?                ��#��@��/����?                ��/����?        ��#��@                ��#���?                z�5��@                �k(��2@                ��#���?                ��,���1@                ,�����;@:l��F:R@��8��8:@,�����;@>��18N@H�4H�4@z�5��@�cp>�9@0#0#@z�5��@��On�(@0#0#@z�5��@�cp>'@                E�JԮD!@        z�5��@�cp>@        z�5��@                        �cp>@                ��/����?                ��/����?                ��/����?0#0#@                0#0#@        ��/����?                ���-��*@                ��/����?                ��On�(@        |�5��8@E�JԮDA@0#0# @��#��0@��/���>@        ��#��0@�cp>7@        ��#��@/����/3@        z�5��@0����/@        z�5��@                        0����/@                �cp>@                ��/����?        ��#���?��|��,@                �cp>'@        ��#���?�cp>@        ��#���?                        �cp>@        |�5��(@��/���@        |�5��(@��/����?        �k(��"@                ��#���?                ��#�� @                z�5��@��/����?                ��/����?        z�5��@                        ��/����?                ��/���@                ��/����?                �cp>@        ��#�� @��/���@0#0# @��#�� @        0#0# @                0#0# @��#�� @                        ��/���@                ��On�(@��+��+4@        ��On�(@H�4H�4(@        ��On�(@0#0# @        �cp>@�C=�C=@                0#0#@        �cp>@H�4H�4@        ��/����?                ��/����?H�4H�4@                0#0# @        ��/����?0#0#�?        ��/����?                        0#0#�?        0����/#@0#0#�?        ��/���@0#0#�?        ��/���@                        0#0#�?        �cp>@                        0#0#@                0#0# @�#���I@鰑5@�C=�C=,@�#���I@���-��@H�4H�4@<��,��D@�cp>@        <��,��4@�cp>@        ��#��0@                ��#��@�cp>@        ��#���?�cp>@        ��#���?                        �cp>@        z�5��@                ��#���?                ��#�� @                <��,��4@                <��,��$@��/����?H�4H�4@<��,��$@��/����?0#0#�?<��,��$@��/����?        �k(��"@                ��#���?��/����?        ��#���?                        ��/����?                        0#0#�?                0#0# @        ��|��,@#0#0&@        D�JԮD!@                �cp>@#0#0&@        �cp>@H�4H�4@        �cp>@0#0#�?        �cp>@                        0#0#�?                ��+��+@                ��+��+@��#���?0����/@S2%S2%1@                �C=�C=@��#���?0����/@��+��+$@        ��/����?        ��#���?��/���@��+��+$@��#���?                        ��/���@��+��+$@        ��/����?                ��/����?��+��+$@        ��/����?H�4H�4@        ��/����?0#0#�?                0#0#�?        ��/����?                        0#0# @                �C=�C=@���>��<@;l��F:B@;�;�V@�k(���5@��/���.@0#0# @�k(���5@��/���.@H�4H�4@<��,��4@/����/#@        �P^Cy/@0����/@                ��/����?        �P^Cy/@��/���@        \Lg1��&@��/����?        ;��,��$@                ��#���?��/����?                ��/����?        ��#���?                ��#��@�cp>@                �cp>@        ��#��@                ;��,��@0����/@        ��#���?��/���@        ��#���?                        ��/���@        ��#��@��/����?        ��#��@                ��#���?                z�5��@                        ��/����?        ��#���?�cp>@H�4H�4@        ��/����?H�4H�4@                H�4H�4@        ��/����?        ��#���?��/���@        ��#���?��/����?                ��/����?        ��#���?                        �cp>@                ��/����?                ��/����?                        ��+��+@                0#0#�?                0#0#@���>��@鰑5@�ڬ�ڬT@���>��@/����/3@�A�A>@z�5��@0����/3@�C=�C=,@��#��@E�JԮD1@H�4H�4@��#��@���-��@��+��+@��#�� @��/����?        ��#�� @                        ��/����?        ��#�� @0����/@��+��+@        �cp>@        ��#�� @��/����?��+��+@��#�� @��/����?0#0# @        ��/����?0#0# @                0#0# @        ��/����?        ��#�� @                                H�4H�4@        鰑%@0#0#�?                0#0#�?        鰑%@        ��#�� @��/����?0#0# @��#���?                ��#���?��/����?0#0# @��#���?��/����?0#0# @        ��/����?0#0# @                ��+��+@        ��/����?H�4H�4@        ��/����?                        H�4H�4@��#���?                        ��/����?        ��#���?        0#0#0@                �C=�C=,@��#���?        0#0# @                0#0# @��#���?                        ��/����?��8��8J@                ��-��-E@        ��/����?��+��+$@        ��/����?                        ��+��+$@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJf��'hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKӅ�h��B(.         �                 ���?��V��O�?)      4�aЁ}@       �                 ��?r?��?�;�?�       ����>u@       �                 0�S�?��p�/_�?�       s0;��r@       �                 @���?���֞F�?�       *�}��r@                          �G�?�V��F
�?�       $�*�q@                        p1�?�=��l�?       <X�a�E@                        ���R?�z�BC��?       �jϦ%�A@                        `&�k?(r��lB�?       ��%��t/@	                        p�x[?���/��?       6��o��#@
                        ���8?��|��?       ���ĺw@                        `7p.?t@ȱ��?       om���S@                        ��>v?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��/���@������������������������       �               ��#���?                        �@�?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �      ��       �cp>@                        ���N?�[nD���?       ���y�O3@                         �!�?��n��?       �-H�\@                        ��y�?�֪u�_�?       ��?�8@������������������������       �               0����/@������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               ��On�(@                        Љ�?��6L�n�?       �E#��h @������������������������       �      �<       ���>��@������������������������       �      ȼ       ��/����?       <                 �&pX?\�:;���?�       ?+D�|\n@        !                 0��?�T`�[k�?.       T��+S@������������������������       �               ��/����?"       5                 pt"?�o;&\��?-       ��e�_�R@#       (                  �f%?��{@��?        )S��aK@$       %                 @*tC?��6L�n�?       ��4}i�8@������������������������       �      �<       �k(���5@&       '                    �?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?)       4                 ��Ɲ?�Z�	7�?       ���`�$>@*       3                 �}kK?��k{��?       _;�W� :@+       .                 �QZ?ذD���?       ������6@,       -                 @F���6L�n�?       �E#��h @������������������������       �      �<       ���>��@������������������������       �      ȼ       ��/����?/       2                 �4Iw?��k*���?       ���b-@0       1                 �L�^?2�c3���?       �uk��!@������������������������       �               0����/@������������������������       �               ��#��@������������������������       �      ȼ       �cp>@������������������������       �               z�5��@������������������������       �               ��#��@6       9                 0��{?�N:�*ط?       I�G�3@7       8                 �m�?      �<       [Lg1��&@������������������������       �               ��#���?������������������������       �               <��,��$@:       ;                 H(�P?x�6L�n�?       �E#��h @������������������������       �               ��/����?������������������������       �      �<       ���>��@=       N                 ���?&�<cgJ�?i       �ͺ���d@>       I                 @+{�?҈�-X�?       s����B@?       @                 �=��?��\���?       �̑-`R9@������������������������       �               ��On�(@A       H                  ���?^�T��?	       ��R�)@B       G                  �/�?� �_rK�?       J�@��"@C       F                 @,G�?�_�A�?       炵�e`@D       E                  ���?�����?       �O��@������������������������       �               ��/����?������������������������       �      �<       ;��,��@������������������������       �      ȼ       ��/����?������������������������       �      �<       ��/����?������������������������       �      ȼ       ��/���@J       K                  y��?����?	       �Ä�>c(@������������������������       �      �<       ���>��@L       M                  �~��?
4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @O       P                 ppla?���+@��?P       �G��f#`@������������������������       �               ��/���@Q       R                 ����?Т�F��?N       �'�5Q_@������������������������       �               ;��,��$@S       f                 @��?�.7iz@�?J       ߉.��\@T       e                 |8��?��r'��?       ``H�#p<@U       Z                  �6�?h�z��P�?       =0F��m;@V       Y                 `U�?)���?       y��uk!@W       X                 x5W�?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �               �cp>@[       `                    �?BG@^���?        X;�8�2@\       ]                 0�M�?���};��?       ��;̑�%@������������������������       �               H�4H�4@^       _                  `���?l�4���?       �tCP��@������������������������       �               �cp>@������������������������       �               0#0# @a       d                 �M��?�@G���?       hu��@b       c                 ���?      �<       �cp>@������������������������       �               ��/����?������������������������       �               0����/@������������������������       �               0#0# @������������������������       �               0#0#�?g       �                  ��^�?��OW�Q�?8       �w4��U@h       w                 \F�M?]����?*       ��'qO@i       t                 `bS�?V�	��`�?       �I9 �1@j       m                 @ۣ?�6�D��?       w�/@k       l                 �#8~?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@n       o                 ���?$I�cͿ�?
       ��J#�l'@������������������������       �               ���-��@p       s                  �g<�?��b�}�?       ���\�@q       r                  $��?X����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �      ��       ��/����?u       v                 ��x�?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?x       �                  �[??2~46�?       !wz��F@y       ~                 Oz�?�,�a�z�?       ��$hB@z       {                 `��?��t� �?       ����x&@������������������������       �               ��#�� @|       }                 �1�?V%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?       �                 `TF�?���~��?       ]����8@������������������������       �      �<       ZLg1��6@�       �                 �C8�?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?�       �                 �;[?tR����?       p\����!@�       �                  �a�?��íxq�?       $2��-�@������������������������       �               �cp>@�       �                 ����?��q�R�?       C}Ԥ@�       �                 P���?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               z�5��@�       �                 `��\?�d��6�?       䰒��7@�       �                 pEʦ?����e�?       �S�)�4@�       �                    �?@ǵ3���?       �q�ͨ�@�       �                 GҎi?��|��?       ���ĺw@������������������������       �               0����/@������������������������       �               ��#�� @������������������������       �               ��#���?�       �                   Y��?*@�����?       \n\�/V)@������������������������       �               D�JԮD!@������������������������       �               0#0#@������������������������       �               H�4H�4@������������������������       �     `=       H�4H�4@�       �                �Y�X�?�=s{Ab�?       aI��n'@������������������������       �               0#0#�?�       �                 �D�1?      �<       鰑%@������������������������       �               ��/���@������������������������       �               ���-��@�       �                 �/O�?Hl���k�?       �-]ƗC@�       �                  ����? L�0�h�?       k�e�C@�       �                 ��_�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                  �!�?Pʊs`�?       �	S\!B@������������������������       �      м       =�C=�C?@�       �                 @��?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?������������������������       �      �<       ��/����?�       �                  �fq?�;�dW��?S       W�;��`@�       �                 `�d�?�(���C�?,       ��a�L6R@�       �                   .p�?�D��7��?       �5�<��F@������������������������       �               ���-��@�       �                 �gY�?��pUз?       }�w�C@�       �                    �?�	6?�?       ���J��A@�       �                 �}��?t��ճC�?       y��l$,@������������������������       �               H�4H�4(@�       �                 �!�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 ���?      �<       ��-��-5@������������������������       �               0#0# @������������������������       �               ��)��)3@�       �                 H~��?~���|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                 P ��?&b)ǡ��?       xJ���:@�       �                 ���?f%@�"�?       ��[�'@������������������������       �               �cp>@�       �                 P�|�?2�c3���?       �uk��!@������������������������       �               �cp>@�       �                 0�C�?^n����?       � ��w<@������������������������       �               z�5��@�       �                 ����?f%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?�       �                 (I��?�Ԏ�>"�?
       ���p*.@�       �                  �Ԧ�?��('���?	       A�+T*@�       �                 �m��?�D#���?       �B�j@������������������������       �               ��#�� @������������������������       �               0#0#@������������������������       �               �C=�C=@������������������������       �      ȼ       ��/����?�       �                 ��c�?���.��?'       C�C���M@������������������������       �      ȼ       �
��
�E@�       �                 `�r�?x�q����?       O�Q*s�/@������������������������       �               ��/����?�       �                 ����?��E�B��?       dߞKC.@�       �                 �-��?|�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               #0#0&@�t�bh�hhK ��h��R�(KK�KK��h �B�  U^Cyc@N��+c@�fm�f�d@�5��P>b@-����m`@@�C=�CO@�5��P>b@��`@��8��8:@�5��P>b@�����]@k�6k�69@�5��P>b@�����]@#0#06@��b:��*@��|��<@0#0#�?z�5��@�a#6�;@0#0#�?;��,��@鰑%@        ;��,��@0����/@        ��#�� @0����/@        ��#���?0����/@        ��#���?��/����?                ��/����?        ��#���?                        ��/���@        ��#���?                z�5��@                ��#���?                ��#�� @                        �cp>@        ��#���?D�JԮD1@0#0#�?��#���?0����/@0#0#�?        0����/@0#0#�?        0����/@                        0#0#�?��#���?                        ��On�(@        ���>��@��/����?        ���>��@                        ��/����?        ��#��`@���|NV@��-��-5@    �M@E�JԮD1@                ��/����?            �M@��/���.@        ��k(/D@��|��,@        �k(���5@�cp>@        �k(���5@                        �cp>@                ��/����?                ��/����?        �k(��2@�cp>'@        ���>��,@�cp>'@        \Lg1��&@�cp>'@        ���>��@��/����?        ���>��@                        ��/����?        ��#��@鰑%@        ��#��@0����/@                0����/@        ��#��@                        �cp>@        z�5��@                ��#��@                �k(��2@��/����?        [Lg1��&@                ��#���?                <��,��$@                ���>��@��/����?                ��/����?        ���>��@                ��Gp_R@�����Q@��-��-5@���>��,@�cp>7@        ;��,��@&jW�v%4@                ��On�(@        ;��,��@��/���@        ;��,��@��/���@        ;��,��@��/����?        ;��,��@��/����?                ��/����?        ;��,��@                        ��/����?                ��/����?                ��/���@        �k(��"@�cp>@        ���>��@                ��#�� @�cp>@                �cp>@        ��#�� @                    �M@y%jW�vH@��-��-5@        ��/���@            �M@�'�xr�F@��-��-5@;��,��$@                5��tSH@�'�xr�F@��-��-5@��#���?On��O0@#0#0&@��#���?On��O0@��+��+$@��#���?��/���@        ��#���?��/����?                ��/����?        ��#���?                        �cp>@                E�JԮD!@��+��+$@        �cp>@0#0# @                H�4H�4@        �cp>@0#0# @        �cp>@                        0#0# @        �cp>@0#0# @        �cp>@                ��/����?                0����/@                        0#0# @                0#0#�?�,����G@��|��<@��+��+$@�GpAF@��/���.@H�4H�4@���>��@0����/#@0#0#�?;��,��@0����/#@0#0#�?z�5��@��/����?                ��/����?        z�5��@                ��#�� @D�JԮD!@0#0#�?        ���-��@        ��#�� @��/����?0#0#�?��#�� @        0#0#�?                0#0#�?��#�� @                        ��/����?        ��#�� @                ��#���?                ��#���?                �k(��B@�cp>@0#0# @��#��@@��/����?0#0#�?�k(��"@��/����?        ��#�� @                ��#���?��/����?        ��#���?                        ��/����?        �,����7@        0#0#�?ZLg1��6@                ��#���?        0#0#�?                0#0#�?��#���?                ��#��@��/���@0#0#�?��#���?��/���@0#0#�?        �cp>@        ��#���?��/����?0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?��#���?                z�5��@                z�5��@���-��*@�C=�C=@z�5��@���-��*@0#0#@z�5��@0����/@        ��#�� @0����/@                0����/@        ��#�� @                ��#���?                        D�JԮD!@0#0#@        D�JԮD!@                        0#0#@                H�4H�4@                H�4H�4@        鰑%@0#0#�?                0#0#�?        鰑%@                ��/���@                ���-��@                �cp>@xb'vb'B@        ��/����?wb'vb'B@        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?eJ�dJ�A@                =�C=�C?@        ��/����?0#0#@                0#0#@        ��/����?                ��/����?        z�5��@鰑5@��8��8Z@z�5��@:l��F:2@I�4H�4H@        E�JԮD!@�z��z�B@        ���-��@                ��/����?�z��z�B@        ��/����?S2%S2%A@        ��/����?��8��8*@                H�4H�4(@        ��/����?0#0#�?        ��/����?                        0#0#�?                ��-��-5@                0#0# @                ��)��)3@        ��/����?H�4H�4@        ��/����?                        H�4H�4@z�5��@/����/#@#0#0&@��#��@��/���@                �cp>@        ��#��@0����/@                �cp>@        ��#��@��/����?        z�5��@                ��#���?��/����?                ��/����?        ��#���?                ��#�� @��/����?#0#0&@��#�� @        #0#0&@��#�� @        0#0#@��#�� @                                0#0#@                �C=�C=@        ��/����?                �cp>@�C=�C=L@                �
��
�E@        �cp>@��8��8*@        ��/����?                ��/����?��8��8*@        ��/����?0#0# @        ��/����?                        0#0# @                #0#0&@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJy"rhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKǅ�h��B�+         <                 �M�y?p$z�>�?#      ��U�ݑ}@       -                 ��]"?bzw��?K       ���`�_@       
                  9U?@9�)\e�?0       :/1_;"T@                        �I?& k�Lj�?	       e*�}#<-@                       �]u?��F���?       :�.�-'@������������������������       �               ��#���?������������������������       �      ��       鰑%@       	                 Ш��?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @                           �?>VBGf��?'       �u�zP@                        �0�?���cE��?       d�coE@                         y��?��+��?       ���|��C@                        ���^?��x_F-�?       x%jW�v8@                        ��B?\����?       �Fx�v�5@                          ��?�N:�*ط?       I�G�3@                        ,*����FO���?       �ߌ$@                        8*��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ��       ��#�� @������������������������       �               �k(��"@������������������������       �      ȼ       ��/����?                        ��?v%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �        	       �P^Cy/@                        $�!�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?                           ��?d�R���?       �\���7@������������������������       �               ���>��@!       ,                  `%+�?Fǵ3���?
       �q�ͨ�/@"       +                 @*tC?��|��?	       ���ĺw+@#       *                 Xy�?4=�%�?       �(J��#@$       %                 �7�<?�`@s'��?       Ei_y,*@������������������������       �               �cp>@&       )                      Ȕfm���?       ��Z�N@'       (                  ���?d%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��/����?������������������������       �               z�5��@������������������������       �      ��       ��/���@������������������������       �               ��#�� @.       ;                 �߯�?8�j���?       �HI�G@/       0                 @��>����X��?       )��֞F@������������������������       �               ��/����?1       6                    �?���+@�?       ���
$F@2       3                 p��v?�	�� ��?       @�x��>@������������������������       �               ���>��<@4       5                �3�q?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?7       :                 0V��?�(߫$��?       0H����*@8       9                 ���E?җZ�	7�?       j~���@������������������������       �               z�5��@������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �      �<       ��/����?=       �                 ��g?r}��9��?�       �_ ��u@>       �                 ��*?��6����?�       �Tg�(�k@?       z                 ���?��jr3�?^       �j��.b@@       a                 p�%h?v�vM��?N       ��О^@A       H                  @?��?��{�Y��?'       ��av{�L@B       C                    �?l7Y���?	       ���r�&@������������������������       �               ��#�� @D       E                 ��ͅ?T����1�?       ��;9�@������������������������       �               ��#���?F       G                  �.�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?I       `                  @���?��+m���?       �%��y&G@J       K                  L��?(�Jg@��?       ��G� �E@������������������������       �               0#0#@L       _                 .��U?l�4���?       �tCP��C@M       P                  �~��?:�,n�?       ���`�B@N       O                 `��}?�;�a
=�?       ��l��@������������������������       �               0#0#�?������������������������       �               �cp>@Q       ^                 �u�?��<X���?       h��Qz>@R       W                 �%�?
�Ϟi�?       ��RE�:@S       T                 @*��?�;[��G�?       �O�;�]!@������������������������       �      ��       �cp>@U       V                   +Y�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?X       ]                  h2�?l����?       �����1@Y       \                 ��}�?z�G���?       ��%�|@Z       [                 ��q�?�@����?       ���a�@������������������������       �               ��/����?������������������������       �               0#0#@������������������������       �               �cp>@������������������������       �               ��+��+$@������������������������       �      м       ��/���@������������������������       �      �<       ��/����?������������������������       �      �<       z�5��@b       o                 p�ʞ?p��x���?'       �!��4P@c       d                     �?h�އQ�?       Շ(�fC@������������������������       �               �cp>@e       l                 �f�?D6��l�?       ���Aj�A@f       i                 @��?0�#�ݬ?       0X{Z�@@g       h                 ��Lx?�����?       �O��@������������������������       �               ��/����?������������������������       �               ;��,��@j       k                 ��
n?      �<       ��b:��:@������������������������       �               ��#�� @������������������������       �               |�5��8@m       n                 P�|�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?p       w                 �ì?�&�K�?       ��l�:@q       v                  0Y��?@n~�ZZ�?
       ���x�U1@r       u                 ���?����?	       !I0`�,@s       t                  ��g�?�FO���?       �ߌ$@������������������������       �               ��/����?������������������������       �               �k(��"@������������������������       �               0#0#@������������������������       �               H�4H�4@x       y                  h��?�;[��G�?       �O�;�]!@������������������������       �      �<       ��/���@������������������������       �               0#0#�?{       �                  �@�?���5r�?       ��#�%�6@|       �                 �_��?��O�:�?       �ʒ�6@}       �                 @�ٿ?��;�� �?       ).���4@~       �                 �L�?B0�8���?
       "Z��!�)@       �                  P�"�?�v�;B��?       ՟���	 @������������������������       �               ��/����?������������������������       �               �C=�C=@�       �                 �D��d�4���?       �tCP��@�       �                 H ȶ?�@G���?       hu��@�       �                 hW�?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               0#0# @������������������������       �      �<       ��#���?������������������������       �      �<       ��/����?�       �                 pb�?ҡ掇��?3       ��5��S@�       �                 \F�M?�M�a���?       |�Pa�qE@�       �                 s��?� N��?       �L�EBC3@������������������������       �               ���-��*@�       �                 `P��?t@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@�       �                    �?jSmd�d�?       -D�|\�7@�       �                 0���?ʔfm���?       ��Z�N/@�       �                 �N�?�`@s'��?
       Ei_y,*+@�       �                 ���s?`n����?       � ��w<@������������������������       �               ��#���?�       �                 (�2�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 p��A?      �<       鰑%@������������������������       �               �cp>@������������������������       �               ��/���@������������������������       �               ��#�� @�       �                 �ؙ�?�̥Q)�?       �9C�<�@�       �                  n��?    ��?       "F�b@������������������������       �               ��#�� @������������������������       �               H�4H�4@������������������������       �      ȼ       �cp>@�       �                 @�C�?4K@�Y{�?       ����A@�       �                 �AS?����|e�?       �z �B�@������������������������       �               ��+��+@�       �                 �C��?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                   E(�?j�\U��?       ]�u��;@�       �                 p��?e��}�?       ��Se+@������������������������       �               ��On�(@������������������������       �      �<       ��#���?�       �                 0�5�?N�;3C(�?
       ��V�s,@�       �                    �?�����?       �O��@������������������������       �               ��/����?������������������������       �               ;��,��@�       �                 XO�?�~�&��?       ?�]��@������������������������       �               ��+��+@������������������������       �               �cp>@�       �                 P���?���Y<'�?G       �Բ��^@�       �                    �?@in��?9       �����X@������������������������       �      ܼ       ������J@�       �                 p?�?.!�4��?       �l���kF@�       �                 @F����J���?        g�챂B@�       �                 X�;�?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?�       �                 8�C�?��i���?       ����A@������������������������       �      ��       %S2%S27@�       �                 ����?�'z�3�?       ���da�%@�       �                 ���?���mf�?       毠�?b@������������������������       �      �<       ��/���@������������������������       �               0#0#�?������������������������       �               H�4H�4@�       �                 �j��?�ǧ\�?       �,W J@������������������������       �      ��       0����/@������������������������       �               H�4H�4@������������������������       �               H�4H�48@�t�bh�hhK ��h��R�(KK�KK��h �B�  	��GPd@E�JԮDa@��N�Ďe@����JW@�-����@@        �#���I@��|��<@        z�5��@�cp>'@        ��#���?鰑%@        ��#���?                        鰑%@        ��#�� @��/����?                ��/����?        ��#�� @                5��tSH@D�JԮD1@        ��,���A@��/���@        ��,���A@0����/@        ������3@0����/@        �k(��2@�cp>@        �k(��2@��/����?        �k(��"@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                �k(��"@                        ��/����?        ��#���?��/����?                ��/����?        ��#���?                �P^Cy/@                        �cp>@                ��/����?                ��/����?        ��b:��*@0����/#@        ���>��@                z�5��@/����/#@        ��#��@0����/#@        ��#��@�cp>@        ��#���?�cp>@                �cp>@        ��#���?�cp>@        ��#���?��/����?        ��#���?                        ��/����?                ��/����?        z�5��@                        ��/���@        ��#�� @                <��,��D@0����/@        =��,��D@��/���@                ��/����?        >��,��D@�cp>@        Jp�}>@��/����?        ���>��<@                ��#���?��/����?                ��/����?        ��#���?                [Lg1��&@��/����?        z�5��@��/����?        z�5��@                        ��/����?        ��#�� @                        ��/����?        j1��tVQ@��F:l$Z@��N�Ďe@j1��tVQ@��h
�W@�A�AN@-�����K@��]�ڕE@%S2%S2G@�>��nK@2����/C@�s?�s?=@��b:��*@�cp>7@��-��-5@;��,��$@        0#0#�?��#�� @                ��#�� @        0#0#�?��#���?                ��#���?        0#0#�?��#���?                                0#0#�?z�5��@�cp>7@��+��+4@        �cp>7@��+��+4@                0#0#@        �cp>7@0#0#0@        鰑5@0#0#0@        �cp>@0#0#�?                0#0#�?        �cp>@                ��/���.@�A�A.@        �cp>'@�A�A.@        ��/���@0#0#�?        �cp>@                ��/����?0#0#�?                0#0#�?        ��/����?                ��/���@�C=�C=,@        ��/���@0#0#@        ��/����?0#0#@        ��/����?                        0#0#@        �cp>@                        ��+��+$@        ��/���@                ��/����?        z�5��@                =��,��D@��/���.@0#0# @���b:@@���-��@                �cp>@        ���b:@@��/���@        ���b:@@��/����?        ;��,��@��/����?                ��/����?        ;��,��@                ��b:��:@                ��#�� @                |�5��8@                        �cp>@                ��/����?                ��/����?        �k(��"@D�JԮD!@0#0# @�k(��"@��/����?�C=�C=@�k(��"@��/����?0#0#@�k(��"@��/����?                ��/����?        �k(��"@                                0#0#@                H�4H�4@        ��/���@0#0#�?        ��/���@                        0#0#�?��#���?0����/@S2%S2%1@��#���?��/���@S2%S2%1@        ��/���@S2%S2%1@        ��/���@vb'vb'"@        ��/����?�C=�C=@        ��/����?                        �C=�C=@        �cp>@0#0# @        �cp>@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?                        0#0#�?                0#0# @��#���?                        ��/����?        ��b:��*@p��F:lI@�C=�C=,@���>��@Pn��O@@H�4H�4@��#���?:l��F:2@                ���-��*@        ��#���?0����/@        ��#���?                        0����/@        z�5��@��|��,@H�4H�4@��#��@�cp>'@        ��#�� @�cp>'@        ��#�� @��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                        鰑%@                �cp>@                ��/���@        ��#�� @                ��#�� @�cp>@H�4H�4@��#�� @        H�4H�4@��#�� @                                H�4H�4@        �cp>@        z�5��@:l��F:2@#0#0&@        ��/����?H�4H�4@                ��+��+@        ��/����?0#0#�?                0#0#�?        ��/����?        z�5��@On��O0@��+��+@��#���?��On�(@                ��On�(@        ��#���?                ;��,��@��/���@��+��+@;��,��@��/����?                ��/����?        ;��,��@                        �cp>@��+��+@                ��+��+@        �cp>@                鰑%@Ϸ|˷�[@        鰑%@��o���U@                ������J@        鰑%@T2%S2%A@        �cp>@=�C=�C?@        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/���@�A�A>@                %S2%S27@        ��/���@�C=�C=@        ��/���@0#0#�?        ��/���@                        0#0#�?                H�4H�4@        0����/@H�4H�4@        0����/@                        H�4H�4@                H�4H�48@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�A�'hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKׅ�h��B/         �                 pK�b?d�~twG�?%      �����p}@       �                  ���?Lqd���?�       &���Qv@       4                 @Ws�?�!� �\�?�       E�C�u@                         @(B�?�Qޔ�?4       �j�b�T@                        �/��? J�����?       g�C���3@������������������������       �               ��#��@                        ���>py8�n�?	       O(�\S'/@������������������������       �               ��#�� @	                       ���8?e��}�?       ��Se+@
                       @u}<9?Ȕfm���?       ��Z�N@                        ��p?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��/����?������������������������       �      ��       0����/#@       '                 ��Н?6v�2�?'       �	u-�VO@       $                 �ڡC?H���'0�?       ��)�F@                        �]t?��6L�n�?       ;�=-�D@                        �y�����k\��?       mG�
 B@                        �Q�?���Ѯ�?       ��GQ&@                        @.��>���/��?       Az$S��@������������������������       �               ��#�� @                          �x�?Δfm���?       ��Z�N@                         �~��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��/����?������������������������       �      �<       ;��,��@������������������������       �      ��       z�5��8@       #                 �{{�?�Z�	7�?       j~���@                            �?�����?       ��X�)B@������������������������       �               ��#���?!       "                 l�Zq?bn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?%       &                 ����?      �<       0����/@������������������������       �               ��/����?������������������������       �               ��/���@(       1                 ��~?F����?       �j�2��0@)       *                 @�ߪ?�!�a6Z�?	       ���t0�'@������������������������       �               �cp>@+       ,                 �؉�?��Ϟi�?       ��ؠ�!@������������������������       �               ��/����?-       .                 �7ڶ?�AP�9��?       i��6��@������������������������       �               0#0#@/       0                 �?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?2       3                 �O@�?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?5       �                   p��?���b��?�       �;o¨�p@6       �                 �I��?�+��?�       �XC1[Kn@7       �                 �"��?Щ�=z��?�       n(A+Im@8       q                 ���x?ФQ��?`       ����[�c@9       p                 `Őq?��҄`-�?E       U�޼:\@:       o                 ��=�?�$��?s�?A       �F�X�Z@;       ^                   ��?�;Xl�?=       ǅ��a�X@<       Y                 ���?�P�j���?&       }�~��P@=       V                  T?�}�v�?"       �@��L@>       A                 p�FK?�j��3��?        �2��ܷK@?       @                  ��?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@B       U                  ��?��u��?       3"~���I@C       T                 pZhv?�ۜ�x�?       ���NO,H@D       I                 P�2?̔fm���?       4�x�А3@E       H                 ���?p�r{��?       e�6� @F       G                 `U�?      �<       ���-��@������������������������       �               ��/���@������������������������       �               �cp>@������������������������       �               ��#���?J       K                 �q�3?h%@�"�?       ��[�'@������������������������       �               ��#�� @L       S                 XBmu?$ k�Lj�?       �q��l}#@M       N                     �?���/��?       V��7�@������������������������       �               ��/����?O       P                 0N�e?`n����?       � ��w<@������������������������       �               ��#���?Q       R                 �9 h?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               ��|��<@������������������������       �      �<       H�4H�4@W       X                 \F�M?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?Z       [                    �?X����1�?       �����x"@������������������������       �               z�5��@\       ]                 (�@�?�J���?       a���@������������������������       �               z�5��@������������������������       �               H�4H�4@_       f                 �΢�Zutee�?       ��@@`       e                 ���?��k*���?       ���b-@a       b                    �?`n����?       � ��w<@������������������������       �               z�5��@c       d                 ��hn?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �      ��       D�JԮD!@g       j                    �?�x�<�?       W&b��q1@h       i                  ��?����X��?       &��֞&@������������������������       �               ;��,��$@������������������������       �      ȼ       ��/����?k       l                 ��;?�����?       �O��@������������������������       �               ��#��@m       n                  ���?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �      ��       �cp>@r                        P�xR?��]O]\�?       ���cG@s       |                 ��.�?d#W�+�?       �W�EaD@t       u                 `U�?�hK)�?       �h��K�B@������������������������       �               �,����7@v       y                 P��;?�(߫$��?       2H����*@w       x                   \��?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?z       {                    �?      �<       ;��,��$@������������������������       �               ��#��@������������������������       �               z�5��@}       ~                 `۶�?z%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?�       �                 ���X?      �<       ���-��@������������������������       �               �cp>@������������������������       �               ��/���@�       �                 ��6�?�b2�ë�?6       z�����R@�       �                 h�B?   �~�?       �ZbQg09@�       �                  @?��?������?       2�<��0@������������������������       �               �cp>@�       �                 G҈n?(�Jg@��?       ��G� �%@������������������������       �               H�4H�4@�       �                  ��?�@G���?       hu��@�       �                 �+��?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      ȼ       0����/@�       �                 �se?      �<	       D�JԮD!@������������������������       �               ��/����?������������������������       �               ���-��@�       �                  �H?3Ԋ�b5�?!       ��o�	�H@�       �                  ��^�?���q���?       �D|+�zA@�       �                  mI�?D�A���?       `�b�79@������������������������       �               ��#�� @�       �                 0�I�?r\{��?       �{�P �0@�       �                    �?���_�?       ���e��#@�       �                 ����?s�T���?       ��e[�&@�       �                 8��?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �      ��       ��#�� @������������������������       �               �cp>@�       �                 `�C?&�b���?       �GXvƒ@�       �                 @��?��ڰ�x�?       �K�f�@������������������������       �               0#0#�?������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?�       �                   ���?����h�?       @��o{#@������������������������       �               0#0# @�       �                 @Ws�?xLU���?       h�ҹ^�@������������������������       �               0#0#�?������������������������       �               ���-��@�       �                 <�Q?��,���?       "C�s��,@�       �                   �G�?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �               0����/@������������������������       �               D�JԮD!@������������������������       �      ��       0#0# @�       �                 �&/�?��+�?       ��؜�_6@������������������������       �               ���>��@������������������������       �        	       �A�A.@�       �                 PAC�?�\�yU�?       ��7�1�#@������������������������       �               ��/����?�       �                    �?�v�;B��?       ՟���	 @�       �                 ��B�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               H�4H�4@�       �                   B�?����)��?@       �r�b\@�       �                 p��{?�w�W��?0       ��!�m�T@�       �                 �@�?����4�?       �#�bh�5@�       �                  ���? �*�'�?       J���ׅ2@�       �                 0�!�?�J�A���?
       3����)@������������������������       �               0#0# @�       �                 Ȑ��?�}/W�?	       �r�.�%@�       �                  �.�?      �<       ���-��@������������������������       �               ��/����?������������������������       �               0����/@������������������������       �               0#0#@������������������������       �      ��       �cp>@������������������������       �               H�4H�4@�       �                 p���?0$OA�?"       P�v��N@������������������������       �        
       S2%S2%1@�       �                 �Z�?��L�`��?       �aMF@������������������������       �               ��/���@�       �                 �O�?4ꌆ��?       ���n�D@������������������������       �               �C=�C=,@�       �                 8�C�?��AA#�?       �>�:@������������������������       �               H�4H�4(@�       �                 ��|�?�j.�d��?	       �I���+@������������������������       �               ��/����?�       �                  \h�?�N�+�?       ����*@������������������������       �               ��/����?�       �                 `���?v=���?       � ��R(@�       �                  D�?�@����?       ���a�@�       �                 ���?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �      ��       H�4H�4@������������������������       �               �C=�C=@������������������������       �      ��       =�C=�C?@�t�bh�hhK ��h��R�(KK�KK��h �B(  C����b@��]�ڕe@���~�gb@C����b@-����/c@��8��8J@C����b@�[<���b@;�;�F@�,����G@�_��e�=@��+��+@���>��@��On�(@        ��#��@                z�5��@��On�(@        ��#�� @                ��#���?��On�(@        ��#���?�cp>@        ��#���?��/����?                ��/����?        ��#���?                        ��/����?                0����/#@        ��k(/D@E�JԮD1@��+��+@�YLg1B@/����/#@        �YLg1B@0����/@        ��#��@@�cp>@        ��#�� @�cp>@        z�5��@�cp>@        ��#�� @                ��#���?�cp>@        ��#���?��/����?                ��/����?        ��#���?                        ��/����?        ;��,��@                z�5��8@                z�5��@��/����?        z�5��@��/����?        ��#���?                ��#�� @��/����?                ��/����?        ��#�� @                        ��/����?                0����/@                ��/����?                ��/���@        ��#��@��/���@��+��+@        ���-��@��+��+@        �cp>@                ��/���@��+��+@        ��/����?                ��/����?��+��+@                0#0#@        ��/����?0#0#�?                0#0#�?        ��/����?        ��#��@��/����?        ��#��@                        ��/����?        �#���Y@2��18^@��+��+D@�5��X@4��18^@k�6k�69@�5��X@5��18^@S2%S2%1@��k(/T@<l��F:R@H�4H�4@�GpAF@3����-O@H�4H�4@�GpAF@P!�ML@H�4H�4@�YLg1B@O!�ML@H�4H�4@��#��0@h
��F@H�4H�4@;��,��$@h
��F@H�4H�4@��#�� @h
��F@H�4H�4@z�5��@��/����?                ��/����?        z�5��@                ;��,��@��]�ڕE@H�4H�4@;��,��@��]�ڕE@        ;��,��@��|��,@        ��#���?���-��@                ���-��@                ��/���@                �cp>@        ��#���?                ��#��@��/���@        ��#�� @                ��#�� @��/���@        ��#�� @��/����?                ��/����?        ��#�� @��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                        �cp>@                ��|��<@                        H�4H�4@��#�� @                ��#���?                ��#���?                z�5��@        H�4H�4@z�5��@                z�5��@        H�4H�4@z�5��@                                H�4H�4@������3@��On�(@        ��#��@鰑%@        ��#��@��/����?        z�5��@                ��#���?��/����?                ��/����?        ��#���?                        D�JԮD!@        �P^Cy/@��/����?        ;��,��$@��/����?        ;��,��$@                        ��/����?        ;��,��@��/����?        ��#��@                ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                        �cp>@        �YLg1B@鰑%@        �YLg1B@��/���@        ��,���A@��/����?        �,����7@                ZLg1��&@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ;��,��$@                ��#��@                z�5��@                ��#���?��/����?                ��/����?        ��#���?                        ���-��@                �cp>@                ��/���@        �P^Cy/@�e�_��G@#0#0&@        &jW�v%4@��+��+@        �cp>'@��+��+@        �cp>@                �cp>@��+��+@                H�4H�4@        �cp>@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @        0����/@                D�JԮD!@                ��/����?                ���-��@        �P^Cy/@�a#6�;@H�4H�4@�P^Cy/@��|��,@��+��+@�P^Cy/@��/���@0#0# @��#�� @                ���>��@��/���@0#0# @��#�� @���-��@0#0#�?��#�� @��/����?0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?        ��#�� @                        �cp>@        ;��,��@��/����?0#0#�?;��,��@        0#0#�?                0#0#�?;��,��@                        ��/����?                ���-��@H�4H�4@                0#0# @        ���-��@0#0#�?                0#0#�?        ���-��@                ���-��*@0#0#�?        0����/@0#0#�?                0#0#�?        0����/@                D�JԮD!@                        0#0# @���>��@        �A�A.@���>��@                                �A�A.@        �cp>@�C=�C=@        ��/����?                ��/����?�C=�C=@        ��/����?0#0#�?                0#0#�?        ��/����?                        H�4H�4@        1����/3@6k�6k�W@        /����/3@R��N��O@        ��On�(@vb'vb'"@        ��On�(@H�4H�4@        ���-��@H�4H�4@                0#0# @        ���-��@0#0#@        ���-��@                ��/����?                0����/@                        0#0#@        �cp>@                        H�4H�4@        ���-��@�;�;K@                S2%S2%1@        ���-��@�z��z�B@        ��/���@                �cp>@�z��z�B@                �C=�C=,@        �cp>@%S2%S27@                H�4H�4(@        �cp>@#0#0&@        ��/����?                ��/����?#0#0&@        ��/����?                ��/����?#0#0&@        ��/����?0#0#@        ��/����?0#0#�?                0#0#�?        ��/����?                        H�4H�4@                �C=�C=@                =�C=�C?@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ���hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK߅�h��B�0         �                 �W�?���|T�?#      N��x��}@       �                 h�b?O��M{�?�       ���]�u@       6                 ��3|?Y��l�?�       ָ�@�r@                          �G�?�:�"�?A       �F����Y@       
                  .�H?.µ*A
�?       ��A抌9@                        p�LP?jP�D�?       �A��P?$@������������������������       �               z�5��@       	                 �㐢?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?                        `&�k?�Tu��?
       ����.@                       ��z�?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��On�(@       %                    �?\������?1       1�g��S@                          D&�?
�U���?!       9ߧ�L@                        �rha?�I��X[�?       �h��G@                        �U���P�؈�w�?       q���S#G@                         �%c?�N,u��?       ��u�=@                          �P�?�Z�	7�?       i~���$@                        ���2?\����?       P	K��@������������������������       �               ��#��@                        4t?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      Լ       �cp>@                         �3��?      �<       ������3@������������������������       �               ��#���?������������������������       �               �k(��2@������������������������       �               ��#��0@������������������������       �      �<       ��/����?!       "                 0p-�?���1n�?       <���4�!@������������������������       �               0����/@#       $                 ��t?�zœ���?       IG���t@������������������������       �               0#0#�?������������������������       �               z�5��@&       '                 $ڗ.?��o��^�?       NjO���5@������������������������       �               �cp>@(       )                  �a�?�e�>�?       n�B��3@������������������������       �               z�5��@*       5                 `�9z?)���?
       T�M��)@+       4                 ���x?�oH2.w�?	       �їD́%@,       3                 �m�M?& k�Lj�?       �q��l}#@-       2                 ֐ɓ?Ȕfm���?       ��Z�N@.       1                ��t��?`n����?       � ��w<@/       0                 �/��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �               0����/@������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��#�� @7       <                 `��?�Aq�\X�?o       ]N��)g@8       9                 P�z�?�֪u�_�?	       � Eowj1@������������������������       �               0����/#@:       ;                 �\ͥ?�ǧ\�?       �,W J@������������������������       �               H�4H�4@������������������������       �               0����/@=       �                 0���?}�A;�?f       C��K�d@>       s                 �"��?�l]N?�?X       O*���a@?       P                 Њ�(?P%��j�?@       ��!�Z@@       C                 ��!?T�־+��?       �I��'3L@A       B                 �e?>ǵ3���?       �q�ͨ�@������������������������       �               z�5��@������������������������       �      ��       0����/@D       O                 �b��?xS%it�?       �;��?H@E       F                �Fq??h�j���?       ���z2@������������������������       �               ��/����?G       L                 � ɒ?h�:V��?       �GP�1@H       K                 ����?�����?       �O��@I       J                 X���?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      ��       z�5��@M       N                 ��d?      �<       [Lg1��&@������������������������       �               ��#��@������������������������       �               ���>��@������������������������       �               Jp�}>@Q       T                ��W�3?�u}�:�?!       t��eI@R       S                 �m۶?��h��?       S�D'�@������������������������       �               0#0# @������������������������       �               ;��,��@U       V                 P�2?\�#���?       �W�%u�E@������������������������       �               ���-��@W       h                 `iև?Ȯ��?       �>`�pB@X       e                 �T��?P�_��?       h�͉V�8@Y       d                  `<��?��Xv#�?       (RҀh�4@Z       a                 PPp�?& k�Lj�?       �q��l}3@[       ^                 �S��?`�i�@M�?       ���wzb0@\       ]                 P.�?      �<	       �cp>'@������������������������       �               ��/����?������������������������       �               鰑%@_       `                 ��s?  k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      ��       ��/���@b       c                  ���?      �<       z�5��@������������������������       �               ��#�� @������������������������       �               ��#���?������������������������       �      �<       ��#���?f       g                    �?      �<       ��#��@������������������������       �               ��#�� @������������������������       �               ��#�� @i       p                 �ז�?�djH�E�?	       ^�\m�n(@j       m                 ��U�?X�j���?       ���z"@k       l                �3�r?      �<       ���>��@������������������������       �               ;��,��@������������������������       �               ��#�� @n       o                    �?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?q       r                 �I��?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @t       �                  ���?B��P���?       �Is���@@u       v                 �Ս�?��f^�|�?       ��S�^u@@������������������������       �        	       ��On�(@w       �                  �Ѱ?v�b���?       �@cr4@x       y                  pjS�?PO���?       ��o0@������������������������       �               ��#���?z       {                 ���8?����VV�?
       A�R.�.@������������������������       �               0����/#@|       }                    �?�֪u�_�?       ��?�8@������������������������       �               ��/���@~                        ��S�?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                ��Sl�?�3`���?       .�r��@������������������������       �               0#0# @�       �                 Po0�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      �<       ��#���?�       �                 �N��?[�æ��?       ��t7 �:@�       �                 �$I�?Xx�Lg�?
       ��[���4@������������������������       �               �cp>@�       �                 (��?1����?	       �`O��2@������������������������       �               H�4H�4@�       �                  ���?��]ۀ��?       E���O(@�       �                 `Fe�?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 ��h�?`���X��?       Pà4�4"@������������������������       �               0#0# @������������������������       �      �<       ��#���?�       �                 0*��?      �<       �cp>@������������������������       �               �cp>@������������������������       �               �cp>@�       �                  �E�?0 A[>�?"       �%Z��K@�       �                    �?���?�s�?       �7y}��<@�       �                  �ni??{�̡�?	       �0M��1@������������������������       �               ��/����?�       �                 `r�t?��2(&�?       �e4��\.@�       �                 @M^i?b,���O�?       ���/> @������������������������       �               ��#�� @������������������������       �               H�4H�4@������������������������       �               �C=�C=@�       �                 ����?�@G���?	       X��Q'@�       �                 Tw�?��XnP��?       ѭS`oM%@������������������������       �               ���-��@�       �                 `Gg�?|�G���?       ��%�|@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �      ��       �;�;;@�       �                 p��z?"L�)wU�?Q       -�Ӈ�_@�       �                 h��?������?:       �1�u��U@�       �                  <�1?J;���p�?(       �Z>/�M@�       �                 `Ar�?T��I�?       
�fyD@������������������������       �               ��/����?�       �                 ����?\�*f��?       �@w�C@������������������������       �               ��/����?�       �                 �m��?���3_��?       �ȓ�B@�       �                  �~��?�yo�z�?       A"�-V*6@������������������������       �               ��/����?�       �                 H{Q�?���yŷ?       L�j>�45@�       �                   ��?�D�-,�?       �D'ŰO@������������������������       �               ��+��+@������������������������       �               ��#���?������������������������       �               �A�A.@�       �                  `���?:HA��]�?
       ��Ƣ�.@�       �                 �?��d
���?       f�G�N�@�       �                ��ߜ?Ȕfm���?       ��Z�N@�       �                 X���?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               H�4H�4@������������������������       �               0#0# @�       �                 ���?@�r���?       %��k�3@�       �                 ���:?ܜ�x�?       d��إV#@�       �                  �Ԧ�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��/���@�       �                 @�C�?(^�yU�?       ��7�1�#@�       �                 �X��?d�ih�<�?       ��
@������������������������       �               0#0#@�       �                  �^��?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 ����?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?�       �                  @?��?l��ʁ�?       �pY;Z;@�       �                 H�sA?�����?       ��X�)B @�       �                  ��g�?l����?       P	K��@������������������������       �               ��/����?������������������������       �               z�5��@������������������������       �      ȼ       ��/����?�       �                 ���?џ[;��?       �RDm&93@�       �                 x�1e?�cj����?       f�e�JO&@�       �                 h��?X����1�?       �����x"@�       �                 CJ�?     ��?       "F�b@������������������������       �               H�4H�4@������������������������       �               ��#�� @������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �               0#0# @�       �                    �?      �<       ��+��+D@������������������������       �               ��-��-5@������������������������       �               ��)��)3@�t�b�T     h�hhK ��h��R�(KK�KK��h �B�  �b:���c@1����/c@�6k�6�c@�}��a@*����m`@\��[�eQ@��tӹa@2��18^@��8��8:@���b:P@�+Q��B@0#0# @��#�� @D�JԮD1@        ���>��@�cp>@        z�5��@                ��#���?�cp>@                �cp>@        ��#���?                ��#���?��|��,@        ��#���?��/����?        ��#���?                        ��/����?                ��On�(@        -�����K@%jW�v%4@0#0# @\Lg1��F@0����/#@0#0#�?���#8E@0����/@        ���#8E@��/���@        
�#���9@��/���@        z�5��@��/���@        z�5��@��/����?        ��#��@                ��#�� @��/����?                ��/����?        ��#�� @                        �cp>@        ������3@                ��#���?                �k(��2@                ��#��0@                        ��/����?        z�5��@0����/@0#0#�?        0����/@        z�5��@        0#0#�?                0#0#�?z�5��@                <��,��$@鰑%@0#0#�?        �cp>@        <��,��$@��/���@0#0#�?z�5��@                ��#��@��/���@0#0#�?��#�� @��/���@0#0#�?��#�� @��/���@        ��#�� @�cp>@        ��#�� @��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#���?                        0����/@                ��/����?                        0#0#�?��#�� @                ���khS@]�ڕ��T@H�4H�48@        ��|��,@H�4H�4@        0����/#@                0����/@H�4H�4@                H�4H�4@        0����/@        ���khS@F�JԮDQ@��-��-5@B����R@H�)�BM@�C=�C=@�YLg1R@��/���>@0#0#@|�5��H@���-��@        z�5��@0����/@        z�5��@                        0����/@        ����JG@��/����?        ��#��0@��/����?                ��/����?        ��#��0@��/����?        ;��,��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        z�5��@                [Lg1��&@                ��#��@                ���>��@                Jp�}>@                \Lg1��6@�e�_��7@0#0#@;��,��@        0#0# @                0#0# @;��,��@                ��,���1@�e�_��7@0#0# @        ���-��@        ��,���1@E�JԮD1@0#0# @�k(��"@��/���.@        ;��,��@��/���.@        ��#��@��/���.@        ��#���?��/���.@                �cp>'@                ��/����?                鰑%@        ��#���?��/���@        ��#���?                        ��/���@        z�5��@                ��#�� @                ��#���?                ��#���?                ��#��@                ��#�� @                ��#�� @                ��#�� @��/����?0#0# @��#�� @��/����?        ���>��@                ;��,��@                ��#�� @                ��#���?��/����?                ��/����?        ��#���?                        ��/����?0#0# @        ��/����?                        0#0# @z�5��@�a#6�;@H�4H�4@��#�� @�a#6�;@H�4H�4@        ��On�(@        ��#�� @��/���.@H�4H�4@��#���?��|��,@0#0#�?��#���?                        ��|��,@0#0#�?        0����/#@                0����/@0#0#�?        ��/���@                ��/����?0#0#�?        ��/����?                        0#0#�?��#���?��/����?0#0# @                0#0# @��#���?��/����?                ��/����?        ��#���?                ��#���?                ��#�� @鰑%@�C=�C=,@��#�� @0����/@�C=�C=,@        �cp>@        ��#�� @��/����?�C=�C=,@                H�4H�4@��#�� @��/����?0#0# @��#���?��/����?        ��#���?                        ��/����?        ��#���?        0#0# @                0#0# @��#���?                        �cp>@                �cp>@                �cp>@        ��#�� @鰑%@�
��
�E@��#�� @鰑%@0#0#0@��#�� @��/����?��8��8*@        ��/����?        ��#�� @        ��8��8*@��#�� @        H�4H�4@��#�� @                                H�4H�4@                �C=�C=@        D�JԮD!@H�4H�4@        E�JԮD!@0#0# @        ���-��@                ��/����?0#0# @                0#0# @        ��/����?                        0#0#�?                �;�;;@�P^Cy/@h
��6@��
�pV@�P^Cy/@h
��6@Z��Y��H@z�5��@9l��F:2@��)��)C@��#�� @���-��@=�C=�C?@        ��/����?        ��#�� @0����/@=�C=�C?@        ��/����?        ��#�� @��/���@=�C=�C?@��#���?��/����?��+��+4@        ��/����?        ��#���?        ��+��+4@��#���?        ��+��+@                ��+��+@��#���?                                �A�A.@��#���?�cp>@#0#0&@��#���?�cp>@H�4H�4@��#���?�cp>@                �cp>@                ��/����?                ��/����?        ��#���?                                H�4H�4@                0#0# @��#���?�cp>'@�C=�C=@��#���?D�JԮD!@        ��#���?��/����?        ��#���?                        ��/����?                ��/���@                �cp>@�C=�C=@        ��/����?H�4H�4@                0#0#@        ��/����?0#0# @        ��/����?                        0#0# @        ��/����?0#0#�?        ��/����?                        0#0#�?{�5��(@��/���@#0#0&@z�5��@��/����?        z�5��@��/����?                ��/����?        z�5��@                        ��/����?        z�5��@��/����?#0#0&@z�5��@��/����?H�4H�4@z�5��@        H�4H�4@��#�� @        H�4H�4@                H�4H�4@��#�� @                ��#��@                        ��/����?                        0#0# @                ��+��+D@                ��-��-5@                ��)��)3@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJJ��hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK���h��B�)         �                 ��g?3�G�?.      a��7�}@       �                 `V3�?�<*z6�?�       �*�Xw@       t                 �&�?��(���?�       "�4��5t@       _                 0S�r?T�x4S�?�       �	X���o@       T                 �:W>?|ϟ6>�?~       Z��XS�h@       !                 �b'�?P4����?^       :�_<�b@                        �y����D��!�?       ��
���L@                        �"�M?1�Cx@��?       X�k�3@@	                        p��R?2d�1s��?       #�!-�=6@
                        ��w@?���3�?       ���(+�%@������������������������       �               �cp>@                        ���>���/��?       U��7�@������������������������       �               �cp>@                           �?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �               ZLg1��&@                        �G��?��k�L�?       sk��#@                           �?p�r{��?       e�6� @                        �-�?r@ȱ��?       om���S@������������������������       �               ��/���@                        ��F�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��/����?������������������������       �               0#0# @                         p���?0���OT�?       r�>%,�9@                        P� ?����X��?       &��֞&@������������������������       �               z�5��@                        ��u0?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �      �<	       ���>��,@"       =                 �ih�?N_/k��??       a�B֓*W@#       0                 �j��?P�%A5L�?!       '�f�C�H@$       -                 p�x[?�d�$���?       >��#�>@%       &                 ��?����ӱ�?       � sE�.0@������������������������       �               z�5��@'       *                 X�+$?���/��?       6��o��#@(       )                 ~W�>r@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@+       ,                 �U���      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@.       /                  ��?�=�Sο?	       ����,@������������������������       �               ��/����?������������������������       �      ��       ��b:��*@1       2                 @6� ?�KĈ�?       y�Zc�2@������������������������       �               0����/@3       8                 �R�־�)z� ��?       ��\�,@4       5                  ��g�?r@ȱ��?       om���S@������������������������       �               ��/���@6       7                 �2*�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?9       :                 `xNv?��6L�n�?       �E#��h @������������������������       �      �<       z�5��@;       <                 pU�,?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?>       ?                   ��?���q���?       �4�E@������������������������       �               ��#�� @@       M                 ����?��c����?       T���D@A       J                 �@�? &t���?       Ķ���=@B       C                 ���?<��S���?       �v�:@������������������������       �        	       ��/���.@D       G                    �?"Iz�9��?       ��[%@E       F                  �\�?�`@s'��?       Ei_y,*@������������������������       �               ��#���?������������������������       �               �cp>@H       I                   �?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@K       L                  ���?ln����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?N       S                  ��?�Z'Q���?       ���]�6(@O       R                 �k�?r�T���?       ��e[�&@P       Q                 ��?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               0#0#�?������������������������       �               0#0# @U       V                   s��?x�V"�?         5N�[,G@������������������������       �      �<       �cp>7@W       ^                 p�D�?��n��U�?       6�8XyR7@X       [                 �$I�?2��[Q;�?       J��yIg5@Y       Z                 �-�?z�G���?       '5L�`�@������������������������       �               �cp>@������������������������       �               H�4H�4@\       ]                 Э=e?��%�?        ����.@������������������������       �        
       ���>��,@������������������������       �               0#0#�?������������������������       �      м       ��/����?`       e                 ��8�?��6�
�?&       �	�]ڰL@a       d                 �l�}?<9�)\e�?       _���b @b       c                 �|?�����?       �O��@������������������������       �               ��/����?������������������������       �               ;��,��@������������������������       �      м       ��/����?f       s                 P #�?lUM�q��?       ܙݰ�H@g       j                  p%+�?T+z8���?       b�0�5/H@h       i                    �?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?k       l                  bB?�?`�W�?       ��d �/G@������������������������       �      ȼ       ������C@m       r                    �?SH����?       ��ϭ
*@n       q                 �Ts�?��Z�	7�?       i~���@o       p                 0���?`%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �               0#0# @������������������������       �      �<       ��/����?u       �                 ��jm?�;?����?0       M"T�IQ@v       �                  ���?��6��?       �m�S=@w       �                 ���?�<;�`(�?       ��^�6@x       y                 H8��?�\z����?       ���U��1@������������������������       �               0#0#@z       �                  `%+�?�Z�ܙ�?       d����+@{       �                 ��:�?�oH2.w�?
       �їD́%@|                        �i�?�֪u�_�?       ��?�8@}       ~                 @aݨ?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?������������������������       �               �cp>@�       �                 @?4=�%�?       �(J��@�       �                  ���?bn����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               ��/����?�       �                  0Y��?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?�       �                 p	o�?      �<       ��#��@������������������������       �               ��#�� @������������������������       �               ��#�� @������������������������       �               �C=�C=@�       �                 @��?��;�,�?       �T��
D@�       �                 pZ9�?2��1 ��?       �w��<@�       �                 �v��?�dI�Ɲ�?       ɑ�P>z2@�       �                 P�<�?�3`���?       .�r��@�       �                 PM@�?���`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               ��#���?�       �                  `s�?��&���?
       ��G2��,@������������������������       �               ��#���?������������������������       �        	       ���-��*@�       �                 p�ռ?ԟ��X�?       m�n�/$@������������������������       �               0#0# @�       �                      u�T���?       ��e[�& @�       �                 @�C�?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?�       �                 0�j�?z��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?�       �                 0vբ?      �<       �cp>'@������������������������       �               ��/����?������������������������       �               0����/#@�       �                  ���?pm�?       �W��3I@�       �                 �!�?c��Q�A�?       �+q��7@�       �                 �b'�?���ʐ��?	       .�i�Pc/@�       �                 (H?d����?       �����!@������������������������       �      ��       �C=�C=@������������������������       �      �<       ��/����?������������������������       �      ��       ���-��@������������������������       �               ��#�� @�       �                 ����?      �<       ��8��8:@������������������������       �               0#0#�?������������������������       �               k�6k�69@�       �                 @�i?y����?A       @ê\�X@�       �                 ��?طB" �?
       ���<�!*@�       �                 ��,z?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               vb'vb'"@�       �                  �E�?�8M�ҿ?7       02�&�U@�       �                 �bW�?4�
Fq�?       /��C@�       �                    �?*^�yU�?       ��7�1�3@������������������������       �               vb'vb'"@�       �                 �yE�?*�Jg@��?       ��G� �%@������������������������       �               ��+��+@������������������������       �               �cp>@�       �                 x�t?      �<       vb'vb'2@������������������������       �               0#0#�?������������������������       �               S2%S2%1@������������������������       �               G�4H�4H@�t�bh�hhK ��h��R�(KK�KK��h �B�  ���#8e@����-�a@�|˷|d@cCy��d@�]�ڕ�`@fJ�dJ�Q@�b:���c@�]�ڕ�_@�z��z�B@�YLg1b@G��t��V@vb'vb'2@�5��X@鰑U@0#0#0@�YLgqT@P!�ML@H�4H�4(@=��,��D@��|��,@0#0# @��#��0@���-��*@0#0# @�P^Cy/@���-��@        ��#��@���-��@                �cp>@        ��#��@��/���@                �cp>@        ��#��@��/����?        ��#��@                        ��/����?        ZLg1��&@                ��#���?���-��@0#0# @��#���?���-��@        ��#���?0����/@                ��/���@        ��#���?��/����?                ��/����?        ��#���?                        ��/����?                        0#0# @|�5��8@��/����?        ;��,��$@��/����?        z�5��@                ��#��@��/����?                ��/����?        ��#��@                ���>��,@                ��k(/D@鰑E@��+��+$@��#��@@On��O0@        |�5��8@�cp>@        \Lg1��&@0����/@        z�5��@                ;��,��@0����/@        ��#���?0����/@        ��#���?                        0����/@        ��#��@                ��#���?                z�5��@                ��b:��*@��/����?                ��/����?        ��b:��*@                ��#�� @鰑%@                0����/@        ��#�� @�cp>@        ��#���?0����/@                ��/���@        ��#���?��/����?                ��/����?        ��#���?                ���>��@��/����?        z�5��@                ��#���?��/����?                ��/����?        ��#���?                ���>��@�cp>�9@��+��+$@��#�� @                ;��,��@�cp>�9@��+��+$@z�5��@��On�8@0#0#�?��#���?�e�_��7@0#0#�?        ��/���.@        ��#���?D�JԮD!@0#0#�?��#���?�cp>@        ��#���?                        �cp>@                �cp>@0#0#�?                0#0#�?        �cp>@        ��#�� @��/����?        ��#�� @                        ��/����?        ��#�� @��/����?vb'vb'"@��#�� @��/����?0#0#�?��#�� @��/����?                ��/����?        ��#�� @                                0#0#�?                0#0# @���>��,@�a#6�;@0#0#@        �cp>7@        ���>��,@0����/@0#0#@���>��,@�cp>@0#0#@        �cp>@H�4H�4@        �cp>@                        H�4H�4@���>��,@        0#0#�?���>��,@                                0#0#�?        ��/����?        4��tSH@���-��@0#0# @;��,��@�cp>@        ;��,��@��/����?                ��/����?        ;��,��@                        ��/����?        �k(���E@��/���@0#0# @�k(���E@�cp>@0#0# @��#���?��/����?                ��/����?        ��#���?                ���#8E@��/����?0#0# @������C@                z�5��@��/����?0#0# @z�5��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                                0#0# @        ��/����?        ���>��,@����z�A@��)��)3@��#�� @��/���@��8��8*@��#�� @��/���@H�4H�4@��#��@��/���@H�4H�4@                0#0#@��#��@��/���@0#0# @��#�� @��/���@0#0#�?        0����/@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@        ��#�� @�cp>@        ��#�� @��/����?        ��#�� @                        ��/����?                ��/����?        ��#�� @        0#0#�?��#�� @                                0#0#�?��#��@                ��#�� @                ��#�� @                                �C=�C=@z�5��@�a#6�;@H�4H�4@z�5��@Nn��O0@H�4H�4@��#�� @��|��,@0#0# @��#���?��/����?0#0# @        ��/����?0#0# @        ��/����?                        0#0# @��#���?                ��#���?���-��*@        ��#���?                        ���-��*@        ��#��@��/����?0#0#@                0#0# @��#��@��/����?0#0# @��#��@��/����?        ��#��@                        ��/����?                ��/����?0#0# @                0#0# @        ��/����?                �cp>'@                ��/����?                0����/#@        ��#�� @E�JԮD!@B�A�@@��#�� @E�JԮD!@�C=�C=@        E�JԮD!@�C=�C=@        ��/����?�C=�C=@                �C=�C=@        ��/����?                ���-��@        ��#�� @                                ��8��8:@                0#0#�?                k�6k�69@��#�� @��/���@��
�pV@��#�� @��/����?vb'vb'"@��#�� @��/����?        ��#�� @                        ��/����?                        vb'vb'"@        �cp>@��+��+T@        �cp>@0#0#@@        �cp>@�C=�C=,@                vb'vb'"@        �cp>@��+��+@                ��+��+@        �cp>@                        vb'vb'2@                0#0#�?                S2%S2%1@                G�4H�4H@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�U�uhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKӅ�h��B(.         v                 �LW�?�v��8S�?&      ��.�}@       s                  d��?t�� 0�?�       ��s�p@       r                 p�3g?�ɠ5y�?�       N��Ǉn@       c                 ��?̃�����?�       �өg�l@       8                 @F����Y�u�?w       E�݃��f@                        ��?�si��?I       u���'�Y@                        �0l?D]8�a��?&       ��S��K@                        �U����X�Ր��?       ��:�QE@	                        p��R?��k{��?       ^;�W� *@
                        ��??��fm���?       ��Z�N@                         _�
?
4=�%�?       �(J��@������������������������       �               ��#�� @������������������������       �               �cp>@������������������������       �      ȼ       �cp>@������������������������       �               ;��,��@                        ��g^?��^��\�?       H��⋣=@                        �5�P?f%@�"�?       ��[�@������������������������       �               ��/����?                         `�J�?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @                        �;�?�q�Ptܳ?       R�� 5�7@������������������������       �        
       �k(��2@                        �2OV?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?                        Ax�@?      �<       �cp>'@������������������������       �               ��/����?������������������������       �               /����/#@       '                 �?B�1����?#       -j���H@       "                  FS?���ae��?       �2��1@        !                  P�J�?�`@s'��?       Ei_y,*@������������������������       �               ��#���?������������������������       �               �cp>@#       &                 ��|�?ػ��ʫ�?       eX'xj&@$       %                 x��U?�d�$���?       �T�f$@������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?������������������������       �               0#0#�?(       7                 �jU?x��#n�?       x���?@)       .                 p�?�$jʲ��?       ����>@*       +                 ��?`n����?       � ��w<@������������������������       �               ��#���?,       -                 ܙ?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?/       6                  @(B�?��F��^�?       Ҧ (2	;@0       5                 p��!?wT �+��?       ��>Y��@1       2                 ��?�3`���?       .�r��@������������������������       �               0#0# @3       4                  �0��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      �<       鰑5@������������������������       �      �<       ��#���?9       N                 p'v�?|�t���?.       �
B�vS@:       M                  ��g�?�9�6��?       �l�=#[A@;       L                 �2FE?��b���?       ��N�e@@<       I                 �$�?@s��?       ŗ��1�:@=       @                 ���>|�6L�n�?       ��4}i�8@>       ?                 U��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?A       F                 `%�7?����X��?       (��֞6@B       C                 p�־?�N:�*ط?       I�G�3@������������������������       �        	       �P^Cy/@D       E                @>�?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@G       H                 �!�?dn����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?J       K                    �?��G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ؼ       z�5��@������������������������       �      �<       ��/����?O       P                 @�~?\C�#ڹ�?       �m7F��E@������������������������       �               ���>��@Q       R                   ��?���/��?       �[[�.�A@������������������������       �               ��/���@S       X                 �?Pw?�A&w(�?       �]��@@T       U                 �=�q?�����?       �O��(@������������������������       �               ���>��@V       W                 @�:�?�Z�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@Y       ^                 ��N�?4=�%�?       �(J��3@Z       ]                 xغD?p�r{��?       e�6� @[       \                 ��Z�?      �<       ���-��@������������������������       �               ��/����?������������������������       �               0����/@������������������������       �               ��#���?_       `                 _%?��<��?       t=�x�(@������������������������       �      ȼ       ;��,��@a       b                 �D��?��|��?       ���ĺw@������������������������       �               0����/@������������������������       �               ��#�� @d       q                  �p�?��Hw�'�?       �ח�G@e       f                 P��?D.��_G�?       �>�Q,{E@������������������������       �        
       �P^Cy/@g       l                 `iև?��P��?       U��o;@h       k                 `�w?��[����?       Hl�_A@i       j                 P*�_?|�G���?       ��%�|@������������������������       �      �<       ��/����?������������������������       �               0#0# @������������������������       �               �cp>@m       p                �Y�k�? �"J�?       �y3D�4@n       o                 8���?�+��0��?       �h}��$@������������������������       �               ���>��@������������������������       �      ȼ       H�4H�4@������������������������       �               ;��,��$@������������������������       �               0#0#@������������������������       �      ��	       0#0#0@t       u                  ��3�?�/�8���?       "Z��!�)@������������������������       �               ��/���@������������������������       �      ��       vb'vb'"@w       x                   ���?LgG���?�       $�dN��j@������������������������       �               0����/#@y       �                  t0�?^׷��?|       t�4c��i@z       }                  ���?d{����?7       2�בtNW@{       |                  PV��?�,m:��?       ܃���=&@������������������������       �               ��#���?������������������������       �               ��+��+$@~       �                 ����?�����D�?0       ���Y��T@       �                 �I�?7_�dFK�?)       ŷ��FP@�       �                    �?P�H�q�?'       49�L O@�       �                 ���p?�7S��?       #����>@�       �                 �U�,?
�}��	�?       �q�Zz5@�       �                 �-�?�(�>�?       \�(�'@�       �                  ���?t@ȱ��?       nm���S@������������������������       �      ��       0����/@������������������������       �               ��#���?������������������������       �               H�4H�4@�       �                  b9�?      �<       0����/#@������������������������       �               ��/����?������������������������       �               D�JԮD!@������������������������       �               vb'vb'"@�       �                  9ר?�)���?       bO���r?@�       �                 `��?��BG_��?       ���M�U3@������������������������       �               0#0#�?�       �                  �G?�?��%�g�?       ���*wS2@�       �                 ����?�0�~��?       r��GQ1@������������������������       �      ��	       ��On�(@�       �                 ��N�?���mf�?       寠�?b@������������������������       �               0#0#�?������������������������       �      ��       ��/���@������������������������       �               0#0#�?�       �                 `uЭ?s�T���?       Q��z:(@������������������������       �               H�4H�4@�       �                 P3"!?`n����?       ~��Y-"@������������������������       �               ��/����?�       �                  ;ޠ?T����?       P	K��@������������������������       �               ��/����?������������������������       �               z�5��@�       �                  ���?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ��#�� @�       �                  }~�?�Jn�� �?       �+�i�0@������������������������       �               �cp>@������������������������       �               �C=�C=,@�       �                 �2*�?ڀYLy�?E       ���4� \@�       �                 �U��?����A.�?2       ���U
S@�       �                 0�i�?V�d�!L�?        ^�S�9�H@�       �                 0���?�@�܌�?       ��J"y�D@�       �                 `�4x?l�K�+:�?       �ޖ��B@�       �                  R��?vutee�?       �ǟf��8@�       �                 ��w�?�����?       �v�qp�1@�       �                 ��:�?�@����?       ���a�#@������������������������       �               ��+��+@�       �                 Z��?hutee�?       Q9��@�       �                 �/��?����|e�?       �z �B�@�       �                 ����?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               ��/���@������������������������       �               �C=�C=@������������������������       �      ��       ��8��8*@�       �                  �6��?��T���?       ��e[�&@������������������������       �               ��#�� @�       �                 ����?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 �"�?      �<       0#0# @������������������������       �               0#0# @������������������������       �               H�4H�4@������������������������       �               ��8��8:@�       �                  y��?(`S��V�?       LL��L�A@�       �                  V��?r-�E�T�?       ��<)@�       �                 �fC�?�}	;	�?       vK�>4%@������������������������       �               0#0#�?������������������������       �               0����/#@������������������������       �               0#0# @�       �                 ��|�?�1�k(5�?       ��$<7@�       �                 0@�?>�Uzb,�?	       W���bn.@�       �                  Џ~�?�D�-,�?       �D'ŰO@������������������������       �               ��#���?������������������������       �               ��+��+@�       �                  ��?���A���?       ��\�F"@�       �                 ���?l����?       P	K��@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?�       �                 V���?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 ����?w�;B��?       ՟���	 @������������������������       �               �C=�C=@������������������������       �      ȼ       ��/����?�t�bh�hhK ��h��R�(KK�KK��h �B�  g:��,&c@�JԮDmc@�N��Nld@��#��`@��]�ڕU@��)��)C@��#��`@�)�B�T@�s?�s?=@��#��`@�)�B�T@��8��8*@~�5��X@�JԮDmS@0#0#@]Lg1��F@\�v%jWK@H�4H�4@���b:@@h
��6@        ���b:@@鰑%@        ���>��@�cp>@        ��#�� @�cp>@        ��#�� @�cp>@        ��#�� @                        �cp>@                �cp>@        ;��,��@                |�5��8@0����/@        ��#�� @��/���@                ��/����?        ��#�� @��/����?                ��/����?        ��#�� @                \Lg1��6@��/����?        �k(��2@                ��#��@��/����?        ��#��@                        ��/����?                �cp>'@                ��/����?                /����/#@        ��b:��*@Pn��O@@H�4H�4@�k(��"@��/���@0#0#�?��#���?�cp>@        ��#���?                        �cp>@        ��#�� @��/����?0#0#�?��#�� @��/����?        ��#�� @                        ��/����?                        0#0#�?��#��@��On�8@0#0# @z�5��@��On�8@0#0# @��#�� @��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                ��#���?�e�_��7@0#0# @��#���?�cp>@0#0# @��#���?��/����?0#0# @                0#0# @��#���?��/����?                ��/����?        ��#���?                        ��/����?                鰑5@        ��#���?                ��b:��J@�cp>7@0#0#�?*�����;@�cp>@0#0#�?+�����;@��/���@0#0#�?�k(���5@��/���@0#0#�?�k(���5@�cp>@        ��#���?��/����?        ��#���?                        ��/����?        <��,��4@��/����?        �k(��2@��/����?        �P^Cy/@                z�5��@��/����?                ��/����?        z�5��@                ��#�� @��/����?        ��#�� @                        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?z�5��@                        ��/����?        �#���9@E�JԮD1@        ���>��@                �k(��2@E�JԮD1@                ��/���@        �k(��2@���-��*@        ;��,��$@��/����?        ���>��@                z�5��@��/����?                ��/����?        z�5��@                ��#�� @�cp>'@        ��#���?���-��@                ���-��@                ��/����?                0����/@        ��#���?                ���>��@0����/@        ;��,��@                ��#�� @0����/@                0����/@        ��#�� @                ��#��@@0����/@vb'vb'"@��#��@@0����/@��+��+@�P^Cy/@                ��,���1@0����/@��+��+@        0����/@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @        �cp>@        ��,���1@        H�4H�4@���>��@        H�4H�4@���>��@                                H�4H�4@;��,��$@                                0#0#@                0#0#0@        ��/���@vb'vb'"@        ��/���@                        vb'vb'"@;��,��4@E�JԮDQ@D�C=�C_@        0����/#@        <��,��4@�_��e�M@B�C=�C_@[Lg1��&@;l��F:B@;�;�F@��#���?        ��+��+$@��#���?                                ��+��+$@<��,��$@<l��F:B@eJ�dJ�A@<��,��$@�-����@@��-��-5@���>��@�-����@@��-��-5@��#���?��|��,@�A�A.@��#���?��|��,@H�4H�4@��#���?0����/@H�4H�4@��#���?0����/@                0����/@        ��#���?                                H�4H�4@        0����/#@                ��/����?                D�JԮD!@                        vb'vb'"@z�5��@0����/3@H�4H�4@        On��O0@H�4H�4@                0#0#�?        On��O0@0#0# @        On��O0@0#0#�?        ��On�(@                ��/���@0#0#�?                0#0#�?        ��/���@                        0#0#�?z�5��@�cp>@H�4H�4@                H�4H�4@z�5��@�cp>@                ��/����?        z�5��@��/����?                ��/����?        z�5��@                z�5��@                ��#���?                ��#�� @                        �cp>@�C=�C=,@        �cp>@                        �C=�C=,@�k(��"@�cp>7@�6k�6�S@��#�� @鰑%@P��N��O@��#�� @鰑%@�z��z�B@��#�� @鰑%@�s?�s?=@        /����/#@�C=�C=<@        0����/#@�A�A.@        0����/#@0#0# @        ��/����?0#0# @                ��+��+@        ��/����?H�4H�4@        ��/����?H�4H�4@        ��/����?0#0#�?                0#0#�?        ��/����?                        0#0# @        ��/����?                ��/���@                        �C=�C=@                ��8��8*@��#�� @��/����?0#0#�?��#�� @                        ��/����?0#0#�?        ��/����?                        0#0#�?                0#0# @                0#0# @                H�4H�4@                ��8��8:@���>��@��On�(@0#0#0@        0����/#@H�4H�4@        0����/#@0#0#�?                0#0#�?        0����/#@                        0#0# @���>��@�cp>@��8��8*@���>��@��/����?H�4H�4@��#���?        ��+��+@��#���?                                ��+��+@z�5��@��/����?0#0#�?z�5��@��/����?        z�5��@                        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?�C=�C=@                �C=�C=@        ��/����?        �t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJW��]hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK���h��B�5                          `Fe�?%���<�?8      ��i}@                        �Y��?2f辭}�?       9꜊v�@@                        (n�q?pUM�q��?       ڙݰ�8@                        P���>��sx�?       �iۍѧ7@                         ������?       ��X�)B @                         �Q�?��Z�	7�?       j~���@������������������������       �               z�5��@������������������������       �      �<       ��/����?	       
                 h���>      �<       z�5��@������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �      ��       �P^Cy/@������������������������       �               0#0#�?                        �G��?�`���6�?       /u��֝!@                        `��?3y�d��?       �)h�2@                         ���?���mf�?       毠�?b@������������������������       �               �cp>@                        ��ib?~�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?                        �72[?b%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               0#0#�?       �                 p��?�Z��?$      ����Q{@       �                 �8U|?z̒B��?�       ���G�v@       �                   p��?2�|R�?�       �g�6�It@       �                 �&�?���fJ�?�       X�͋^�r@       x                 _5?��|�8�?�       ��?6�l@       3                 ��k?���]��?f       D�zU)<b@       *                 `<��?lQ��?       ��Я[[:@        )                  �0��?)���?       y��uk1@!       (                    �?��i�@M�?       ���wzb0@"       %                 �.��?�F���?       ;�.�-'@#       $                 @�Z�>      �<       D�JԮD!@������������������������       �               ��/����?������������������������       �               ��/���@&       '                 X��?^%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               0����/@������������������������       �      �<       ��#���?+       ,                 @vn?8�c3���?       �uk��!@������������������������       �               z�5��@-       2                 p�e?r@ȱ��?       nm���S@.       /                 �.��?\%@�"�?       ��[�@������������������������       �               ��/����?0       1                  Џ~�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               �cp>@4       W                 0�ӎ?(�0�B�?S       -G�{�]@5       @                  [�f?(�6N�?*       ��ʲ�!M@6       9                  ����?�(߫$��?       3H����:@7       8                 �a?��Z�	7�?       j~���@������������������������       �      �<       z�5��@������������������������       �      ��       ��/����?:       =                 йϷ?�:�^���?       ��]�ڕ5@;       <                 ����?      �<       �k(��2@������������������������       �               ��#���?������������������������       �               ��,���1@>       ?                  ��z?b%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?A       T                 �;�?�-��؈�?       ps�vB�?@B       O                  �!�?��U�ho�?       �wb���;@C       L                 ��ͅ?͏BC��?       �WDl��0@D       G                 wu?x�����?	       �4^$4�#@E       F                 �B{|?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @H       I                 ����?�`@s'��?       Di_y,*@������������������������       �               ��/���@J       K                 hl��?^%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?M       N                 X��?�Qk��?       ��Th!�@������������������������       �               �cp>@������������������������       �               0#0#@P       Q                 ��N�?8k�"O��?       �?<��*&@������������������������       �      �<       z�5��@R       S                  '�?  k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      ��       ��/���@U       V                   ��?      �<       ��/���@������������������������       �               ��/����?������������������������       �               ��/����?X       ]                  `s�? sPVv��?)       ��7�W�N@Y       \                 �=�?$ k�Lj�?       �q��l}@Z       [                �3̳�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               �cp>@^       w                ���ms?�nߡ� �?&       XBe+�1L@_       v                 �$I�?���2�?       '�����@@`       s                  ��?�l��2�?       `���^:@a       b                  h��?��/�{�?        ����:6@������������������������       �               0#0# @c       n                  ����?2��S%�?       �1�F�64@d       e                 )�`f?As.�ʴ�?	        E&A3*@������������������������       �               z�5��@f       g                 #/��?l��w��?       ���@������������������������       �               ��/����?h       k                  @��?��`i��?       �؛.�@i       j                 P]ڒ?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?l       m                 ���?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @o       p                  DŦ?��3Fi�?       :�"Ξs@������������������������       �               H�4H�4@q       r                  `s�?�J���?       ��*]Y@������������������������       �               0#0# @������������������������       �               ��#�� @t       u                 p���?      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@������������������������       �               ���>��@������������������������       �               \Lg1��6@y       �                   s��?<ƙ.U�?9       ��X�U@z       �                  `�J�?�����?       ��9�J5I@{       |                 0�?Zn����?       ~��Y-"@������������������������       �               ��/����?}       ~                    �?T����?       P	K��@������������������������       �               ;��,��@       �                 ����?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                  �e?���P+�?       n�vc��D@�       �                 ���m?)���?       y��uk!@������������������������       �               ��/���@������������������������       �               ��#���?������������������������       �               Qn��O@@�       �                  ��?&����~�?       �rw���@@�       �                 h�B?>�Z���?       _֎V��=@�       �                 ����?��k*���?
       ���b-@�       �                 �Us9?���/��?       U��7�@�       �                 0N?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@�       �                    �?����?       ��X�)B@������������������������       �               ��#�� @�       �                ��3(�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       ���-��@�       �                 �x�?�p����?       �u	h0.@�       �                 `��^?���`�?       ��
�Me@�       �                 �i�?�֪u�_�?       ��?�8@������������������������       �               0����/@������������������������       �               0#0#�?�       �                   �?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               ���>��@�       �                 d�ѣ?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                 �&��?$k�YI��?.        ��P@�       �                  �x��?X�e����?-       �(���P@�       �                 ��?��߁^�?       ��f��>@�       �                 8��?^V�\Ga�?	       q�6t%@�       �                 �^Ҧ?\%��̫�?       �@�o#@������������������������       �               ��#���?�       �                   ҏ�?�;[��G�?       �O�;�]!@�       �                 ��jm?�@G���?       hu��@�       �                 ���?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               ��/����?������������������������       �               0����/@������������������������       �               0#0#�?�       �                �I�s?      �<       %jW�v%4@������������������������       �               �cp>@������������������������       �        
       ��|��,@�       �                 P?��=��?       �֝[:�A@�       �                    �?�4O��?       ���]��9@�       �                 �am�?d�r{��?       e�6� @�       �                  *}�?f%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �               0����/@�       �                 @��?T�b���?       �^Pb
2@�       �                 ����?�]
���?	       ��Ј�'@�       �                 ��ť?޾�R���?       ;�S) $@�       �                  �?��]ۀ��?       E���O@�       �                 p5W�?�@����?       ���a�@�       �                   ���?z��`p��?       �����@������������������������       �               0#0#�?�       �                  `<��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               0#0# @������������������������       �               ��#���?������������������������       �               0#0#@������������������������       �      ȼ       ��/����?�       �                 �n{@?Zn����?       � ��w<@������������������������       �               ��#��@������������������������       �      �<       ��/����?�       �                ��2yt?      �<       /����/#@������������������������       �               0����/@������������������������       �               0����/@������������������������       �     ��<       0#0#�?�       �                 <��?��pI��?       #���D;@�       �                 ��y�?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@�       �                 ��~?FH�=��?       �є�T+6@�       �                  b��>��b�}�?       ���\�@������������������������       �               ��/����?�       �                  @���?T����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @�       �                  ����?,N=� �?       ��a��+1@������������������������       �               0#0#0@������������������������       �      �<       ��#���?������������������������       �     ��       �ڬ�ڬD@�       �                 p��z?�]��t��?.       �G��Q@�       �                 P���?�9}ǀ�?       ���?��:@�       �                 ��?�8f���?       ב+XW�+@�       �                ����}?l@ȱ��?       nm���S@������������������������       �               ��#���?������������������������       �      ��       0����/@�       �                 h��?�~�&��?       ?�]��@�       �                 ��;o?�@����?       ���a�@������������������������       �               H�4H�4@�       �                 ���?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                  �JV�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 pTF�?�n���k�?
       3��&�*@�       �                    �?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               #0#0&@�       �                 ��|�?��К���?       l�[��)F@�       �                 Tw�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                  �?      �<       ��+��+D@������������������������       �               0#0# @������������������������       �               ��)��)C@�t�bh�hhK ��h��R�(KK�KK��h �B�  ��tӹa@��~Y/f@�i��b@[Lg1��6@��/���@H�4H�4@�k(���5@��/����?0#0#�?�k(���5@��/����?        z�5��@��/����?        z�5��@��/����?        z�5��@                        ��/����?        z�5��@                ��#���?                ��#�� @                �P^Cy/@                                0#0#�?��#���?�cp>@0#0# @��#���?�cp>@0#0#�?        ��/���@0#0#�?        �cp>@                ��/����?0#0#�?        ��/����?                        0#0#�?��#���?��/����?        ��#���?                        ��/����?                        0#0#�?+���>�]@����9e@�4H�4�b@    �]@C:l��d@��o���U@    �]@F:l��d@(S2%S2G@
��G�[@������c@�s?�s?=@�#���Y@�B�)[@vb'vb'2@bCy��T@{%jW�vH@��8��8*@z�5��@&jW�v%4@        ��#�� @��/���.@        ��#���?��/���.@        ��#���?鰑%@                D�JԮD!@                ��/����?                ��/���@        ��#���?��/����?        ��#���?                        ��/����?                0����/@        ��#���?                ��#��@0����/@        z�5��@                ��#���?0����/@        ��#���?��/����?                ��/����?        ��#���?��/����?        ��#���?                        ��/����?                �cp>@        ���khS@��|��<@��8��8*@��#��@@鰑5@0#0#@[Lg1��6@��/���@        z�5��@��/����?        z�5��@                        ��/����?        ������3@��/����?        �k(��2@                ��#���?                ��,���1@                ��#���?��/����?        ��#���?                        ��/����?        ;��,��$@E�JԮD1@0#0#@;��,��$@���-��*@0#0#@z�5��@0����/#@0#0#@z�5��@���-��@        ��#�� @��/����?                ��/����?        ��#�� @                ��#���?�cp>@                ��/���@        ��#���?��/����?        ��#���?                        ��/����?                �cp>@0#0#@        �cp>@                        0#0#@���>��@��/���@        z�5��@                ��#���?��/���@        ��#���?                        ��/���@                ��/���@                ��/����?                ��/����?        �GpAF@��/���@vb'vb'"@��#���?��/���@        ��#���?��/����?                ��/����?        ��#���?                        �cp>@        �k(���E@��/���@vb'vb'"@<��,��4@��/���@vb'vb'"@��b:��*@��/���@vb'vb'"@�k(��"@��/���@vb'vb'"@                0#0# @�k(��"@��/���@�C=�C=@���>��@��/���@0#0# @z�5��@                ��#���?��/���@0#0# @        ��/����?        ��#���?��/����?0#0# @��#���?��/����?                ��/����?        ��#���?                        ��/����?0#0# @        ��/����?                        0#0# @��#�� @        ��+��+@                H�4H�4@��#�� @        0#0# @                0#0# @��#�� @                ��#��@                ��#���?                z�5��@                ���>��@                \Lg1��6@                ������3@�_��e�M@��+��+@���>��@��]�ڕE@        z�5��@�cp>@                ��/����?        z�5��@��/����?        ;��,��@                ��#���?��/����?                ��/����?        ��#���?                ��#���?&jW�v%D@        ��#���?��/���@                ��/���@        ��#���?                        Qn��O@@        {�5��(@Nn��O0@��+��+@|�5��(@��/���.@0#0# @��#��@鰑%@        ��#��@��/���@        ��#���?�cp>@        ��#���?                        �cp>@        z�5��@��/����?        ��#�� @                ��#���?��/����?                ��/����?        ��#���?                        ���-��@        ��#�� @0����/@0#0# @��#���?0����/@0#0# @        0����/@0#0#�?        0����/@                        0#0#�?��#���?        0#0#�?��#���?                                0#0#�?���>��@                        ��/����?H�4H�4@        ��/����?                        H�4H�4@���>��@y%jW�vH@#0#0&@���>��@y%jW�vH@��+��+$@��#���?�a#6�;@0#0# @��#���?��/���@0#0# @��#���?��/���@0#0#�?��#���?                        ��/���@0#0#�?        �cp>@0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                ��/����?                0����/@                        0#0#�?        %jW�v%4@                �cp>@                ��|��,@        z�5��@鰑5@0#0# @z�5��@�cp>'@0#0# @��#���?���-��@        ��#���?��/����?                ��/����?        ��#���?                        0����/@        ;��,��@0����/@0#0# @��#���?�cp>@0#0# @��#���?��/����?0#0# @��#���?��/����?0#0#@        ��/����?0#0#@        ��/����?0#0# @                0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?                0#0# @��#���?                                0#0#@        ��/����?        ��#��@��/����?        ��#��@                        ��/����?                /����/#@                0����/@                0����/@                        0#0#�?���>��@�cp>@S2%S2%1@��#��@��/����?                ��/����?        ��#��@                z�5��@��/����?S2%S2%1@��#�� @��/����?0#0#�?        ��/����?        ��#�� @        0#0#�?                0#0#�?��#�� @                ��#���?        0#0#0@                0#0#0@��#���?                                �ڬ�ڬD@��#���?0����/#@!�A�AN@��#���?D�JԮD!@S2%S2%1@��#���?��/���@��+��+@��#���?0����/@        ��#���?                        0����/@                �cp>@��+��+@        ��/����?0#0#@                H�4H�4@        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                ��/����?H�4H�4(@        ��/����?0#0#�?                0#0#�?        ��/����?                        #0#0&@        ��/����?�
��
�E@        ��/����?H�4H�4@        ��/����?                        H�4H�4@                ��+��+D@                0#0# @                ��)��)C@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJt�mUhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK녔h��Bh3         �                 pK�b?��<�P�?(      �;�L{�}@       �                 ���?\(�O��?�       ��{�Vv@       H                 ���?]���Ĩ�?�       �>��&&v@       ;                 ��??L��7�?Z       ����c�a@       ,                 �U����ܘ���?D       ���dcS\@       )                 @G#~?8cpp�R�?(       j}��v�M@                        `f�?&=�U(�?"       ����:�I@                        0�!�?.k�"O��?       �?<��*&@	       
                  P���?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?                         �.�?\����?       P	K��@������������������������       �               ��/����?������������������������       �               z�5��@       "                 wu?l9��;3�?       �ll�D@                         `��?�4��v�?       �Y-"�7@                         ���?��Z�	7�?       ���`�$.@                        ��-�?��k{��?
       _;�W� *@                         ����?@ǵ3���?       �q�ͨ�@������������������������       �               ��#�� @                        @��R?l@ȱ��?       nm���S@������������������������       �      ��       0����/@������������������������       �               ��#���?                         ����?�d�$���?       �T�f@                        ���T?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       z�5��@������������������������       �               ��#�� @       !                    �?)���?       y��uk!@                         �/��?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �               �cp>@#       (                 @��?�O���?
       ��o0@$       '                 Z�K?�Tu��?	       ����.@%       &                 �D�?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �      ��       ��On�(@������������������������       �               0#0#�?*       +                 @���?��6L�n�?       �E#��h @������������������������       �      �<       ���>��@������������������������       �      ȼ       ��/����?-       8                 �c=d?�
O�:��?       ��<�O�J@.       7                 P^N<?���/4��?       ��ƪ�oD@/       0                 �j[?X���m>�?       0w��e�B@������������������������       �               ��b:��*@1       2                 ����?�����?       �O��8@������������������������       �        
       ������3@3       4                 -��?  k�Lj�?       �q��l}@������������������������       �               ��/����?5       6                    �?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      �       �cp>@9       :                 �[V�?   ���?       +x�1�)@������������������������       �               z�5��@������������������������       �      ��       ���-��@<       C                 p��?����β�?       ��D�=;@=       @                  �X?HH�,.̷?       �J�$r.5@>       ?                    �?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?A       B                 �5��>      �<       E�JԮD1@������������������������       �               ��/����?������������������������       �               ��/���.@D       E                 `�??`n����?       � ��w<@������������������������       �               z�5��@F       G                  {X%?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?I       �                  ����?熉5���?�       U��A�j@J       q                 pTF�?��95��?S       h����`@K       L                  ;��?Df�`'��?!       s�B�uK@������������������������       �               z�5��@M       `                 ��*?��8��?       a���ZH@N       U                 u3�?�G���D�?       ���=@O       P                 �aM?�o����?       ���5u*@������������������������       �               ��/����?Q       R                  ����?����X��?       &��֞&@������������������������       �               ��#�� @S       T                  ���?Nn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @V       ]                 ���?�~�&��?	       >�]��/@W       Z                    �?��[����?       Hl�_A@X       Y                 ���?���mf�?       毠�?b@������������������������       �      �<       ��/���@������������������������       �               0#0#�?[       \                 ��9�?v�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?^       _                 �R��?l*�'=P�?        �2"@������������������������       �               0#0# @������������������������       �      ȼ       ��/����?a       b                 0p�:?��t?��?       "���5�3@������������������������       �               0����/@c       h                 ����?rb���?       ���{�-@d       e                 �~�?���WW�?       �j�S@������������������������       �               ��/����?f       g                 |1Ҙ?�|2N��?       �3K}@������������������������       �               z�5��@������������������������       �               0#0# @i       l                  @mj�?����e��?       �ga��!@j       k                  ���?      �<       �cp>@������������������������       �               ��/����?������������������������       �               0����/@m       p                 �Z�?��q�R�?       C}Ԥ@n       o                �Y���?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��#���?r       }                   �G�?^��E�?2       Je��E8T@s       |                 И"�?��|��?       ���ĺw+@t       u                 ����?���/��?       V��7�@������������������������       �               z�5��@v       y                    �?& k�Lj�?       �q��l}@w       x                8�|�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?z       {                 8A!�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �      ��       �cp>@~       �                 0�q�?�P�>���?'       S��`N�P@       �                 ��I�?:S�+�Q�?       �apcc�F@�       �                  ��?�����J�?       P#j|�PE@�       �                 p&͚?)�>�
�?       ����?@�       �                 p`�?\n����?       � ��w<(@�       �                 ��Ӊ?�d�$���?       �T�f$@�       �                 �L�?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ��       ���>��@������������������������       �      ȼ       ��/����?�       �                  @?��?��Z��?       >�mKߣ3@�       �                 |�Յ?L� P?)�?       ����x�@������������������������       �               ��#��@������������������������       �               0#0#�?������������������������       �      ��       ���>��,@�       �                 �ؐ?�it�R��?       ��ǿ%@�       �                     �?���`�?       ��
�Me@������������������������       �               ��#���?�       �                 u�?��[����?       Hl�_A@������������������������       �               0����/@������������������������       �               0#0# @������������������������       �               H�4H�4@������������������������       �      �       �cp>@�       �                 p�Ǩ? c��q��?       �Y�r�5@������������������������       �      ȼ       �P^Cy/@�       �                 `�C?�djH�E�?       ^�\m�n@�       �                 HFU�?L� P?)�?       ����x�@������������������������       �               ��#�� @�       �                 `�>?T����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?�       �                 @aA�?��[����?-       �!�(łS@�       �                 �F��?����(�?$       vo��L�P@�       �                 J�?bn����?       � ��w<8@������������������������       �               ��#��@�       �                 0�!�?�Z�	7�?       j~���4@������������������������       �               �cp>@�       �                 @Ws�?�M:���?	       ����71@������������������������       �      ��       ;��,��$@�       �                  �Mm�?��|��?       ���ĺw@������������������������       �               ��#�� @������������������������       �      ��       0����/@�       �                 ,G�?�Y�����?       ���o]E@������������������������       �               ��+��+$@�       �                 @8x�?,��V�"�?       ��y���?@�       �                 �V�?b�F����?       يj���8@�       �                 ���o?)��G��?       `�o�f�%@������������������������       �               H�4H�4@�       �                 ����?d�r{��?       e�6� @������������������������       �               ��#���?�       �                    �?      �<       ���-��@������������������������       �               0����/@������������������������       �               ��/����?�       �                  ���?�nl4�/�?       SBe+�1,@�       �                �o|?�n���k�?       3��&�*@������������������������       �               vb'vb'"@�       �                 �p�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �      ܼ       ��#���?������������������������       �               �C=�C=@�       �                 0H0�?B������?	       ��Iē'@�       �                 ����?���/��?       Az$S��@������������������������       �               ��/����?�       �                  �E�?�����?       ��X�)B@�       �                 |�y�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                    �?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?�       �                 @  �?�֪u�_�?       ��?�8@������������������������       �               ��/���@�       �                  0Y��?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      �       H�4H�4@�       �                  ����?���q��?L       �O�,��\@�       �                 0�?���OP�?       &��=@�       �                   ��?��[����?       Hl�_A+@������������������������       �               0#0# @�       �                 (��?�֪u�_�?       ��?�8'@�       �                  �?�}	;	�?       vK�>4%@�       �                ���?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               E�JԮD!@������������������������       �               0#0#�?�       �                 �o\�?r����?	       Qz�i0@�       �                 �⊴?|��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �      ��       ��8��8*@�       �                    �?�!����?;       ��E��aU@�       �                   ��?      �<       #0#0F@������������������������       �               0#0#�?������������������������       �               �
��
�E@�       �                   B�?���� ��?       tx[f��D@�       �                 �ڡs?�w��Z��?       �R9@�       �                 ���?h�4���?       �tCP��@������������������������       �               �cp>@������������������������       �               0#0# @�       �                 ����?`,�#6?�?       ���*4@������������������������       �               S2%S2%1@�       �                 |��?���`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      ��       0#0#0@�t�b�!     h�hhK ��h��R�(KK�KK��h �B  ?��,��d@��e�_�b@��
���c@?��,��d@�-����`@�[��[�L@?��,��d@�-����`@�;�;K@������Q@��t�HQ@0#0#�?��#��P@�cp>G@0#0#�?�#���9@On��O@@0#0#�?�k(��2@�]�ڕ�?@0#0#�?���>��@��/���@        ��#���?�cp>@                �cp>@        ��#���?                z�5��@��/����?                ��/����?        z�5��@                [Lg1��&@�a#6�;@0#0#�?;��,��$@���-��*@        �k(��"@�cp>@        ���>��@�cp>@        z�5��@0����/@        ��#�� @                ��#���?0����/@                0����/@        ��#���?                ��#��@��/����?        ��#���?��/����?                ��/����?        ��#���?                z�5��@                ��#�� @                ��#���?��/���@        ��#���?��/����?                ��/����?        ��#���?                        �cp>@        ��#���?��|��,@0#0#�?��#���?��|��,@        ��#���?��/����?                ��/����?        ��#���?                        ��On�(@                        0#0#�?���>��@��/����?        ���>��@                        ��/����?        ��k(/D@���-��*@        Ey�5A@���-��@        Ey�5A@��/���@        ��b:��*@                ;��,��4@��/���@        ������3@                ��#���?��/���@                ��/����?        ��#���?��/����?        ��#���?                        ��/����?                �cp>@        z�5��@���-��@        z�5��@                        ���-��@        ;��,��@h
��6@        ��#���?%jW�v%4@        ��#���?�cp>@                �cp>@        ��#���?                        E�JԮD1@                ��/����?                ��/���.@        ��#��@��/����?        z�5��@                ��#���?��/����?        ��#���?                        ��/����?        �t�Y�W@���|�P@������J@�YLg1R@��]�ڕE@��+��+4@<��,��4@鰑5@��8��8*@z�5��@                ���>��,@鰑5@��8��8*@;��,��$@E�JԮD!@��+��+$@<��,��$@�cp>@                ��/����?        <��,��$@��/����?        ��#�� @                ��#�� @��/����?                ��/����?        ��#�� @                        �cp>@��+��+$@        0����/@0#0# @        ��/���@0#0#�?        ��/���@                        0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?0#0# @                0#0# @        ��/����?        ��#��@��On�(@H�4H�4@        0����/@        ��#��@��/���@H�4H�4@z�5��@��/����?0#0# @        ��/����?        z�5��@        0#0# @z�5��@                                0#0# @��#���?���-��@0#0#�?        �cp>@                ��/����?                0����/@        ��#���?��/����?0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?��#���?                �#���I@h
��6@�C=�C=@��#��@0����/#@        ��#��@��/���@        z�5��@                ��#���?��/���@        ��#���?��/����?                ��/����?        ��#���?                        �cp>@                ��/����?                ��/����?                �cp>@        �,����G@��On�(@�C=�C=@*�����;@�cp>'@H�4H�4@*�����;@D�JԮD!@H�4H�4@��b:��:@��/���@0#0#�?��#�� @��/���@        ��#�� @��/����?        ��#���?��/����?        ��#���?                        ��/����?        ���>��@                        ��/����?        �k(��2@        0#0#�?��#��@        0#0#�?��#��@                                0#0#�?���>��,@                ��#���?0����/@��+��+@��#���?0����/@0#0# @��#���?                        0����/@0#0# @        0����/@                        0#0# @                H�4H�4@        �cp>@        ������3@��/����?0#0#�?�P^Cy/@                ��#��@��/����?0#0#�?��#��@        0#0#�?��#�� @                ��#�� @        0#0#�?                0#0#�?��#�� @                        ��/����?        �k(���5@�cp>7@B�A�@@�k(��2@��/���.@0#0#@@��#��0@��/���@        ��#��@                z�5��(@��/���@                �cp>@        z�5��(@0����/@        ;��,��$@                ��#�� @0����/@        ��#�� @                        0����/@        ��#�� @��/���@0#0#@@                ��+��+$@��#�� @��/���@#0#06@��#�� @��/���@�A�A.@��#���?���-��@H�4H�4@                H�4H�4@��#���?���-��@        ��#���?                        ���-��@                0����/@                ��/����?        ��#���?��/����?H�4H�4(@        ��/����?H�4H�4(@                vb'vb'"@        ��/����?H�4H�4@        ��/����?                        H�4H�4@��#���?                                �C=�C=@z�5��@��/���@0#0#�?z�5��@�cp>@                ��/����?        z�5��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                ��#���?                ��#���?                        0����/@0#0#�?        ��/���@                ��/����?0#0#�?        ��/����?                        0#0#�?                H�4H�4@        ��|��,@s�6k�6Y@        鰑%@��)��)3@        0����/#@0#0#@                0#0# @        0����/#@0#0# @        0����/#@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        E�JԮD!@                        0#0#�?        ��/����?�A�A.@        ��/����?0#0# @                0#0# @        ��/����?                        ��8��8*@        ��/���@�N��NlT@                #0#0F@                0#0#�?                �
��
�E@        ��/���@�z��z�B@        ��/���@��-��-5@        �cp>@0#0# @        �cp>@                        0#0# @        ��/����?��)��)3@                S2%S2%1@        ��/����?0#0# @        ��/����?                        0#0# @                0#0#0@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJc��hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK녔h��Bh3         �                 /O�?^w��K�?+      ���}@       �                 ��g?����?�       �+'�Dv@       �                 0G?�.v~���?�       ��� s@       w                 pTF�?Q��*�?�       �{�̂�o@       l                 �^#�?�[���u�?�       u��wy�k@                        ���a?P>e;��?�       �x���i@                        `���>����ݱ�?       ��"c�ZB@������������������������       �               ��#��@	       
                 �@�F?���3�?       q��^�H@@������������������������       �               z�5��@                        `�yS?jQ��?       ��Я[[:@                        ��g�?������?       �N0gX1@                        @���>Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?                           �?      �<       ���-��*@������������������������       �               ��/����?������������������������       �               ��On�(@                        ��C�?� �_rK�?       J�@��"@                           �?�����?       �O��@                         s��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#��@������������������������       �               �cp>@       %                  L��?H .mK��?m       *�D�YFe@       "                 ���@? =켴��?       �����E@                          ���?x�s�	�?       �rD@                        p�z?p�+�*�?       xȚ�
A@������������������������       �               ��#��@@������������������������       �      �<       ��/����?        !                  `%+�?dn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#��@#       $                 pR��?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?&       9                 `��~?:,?v'�?Q       H�o`@'       (                  h��?$<rW�?       |��z K@������������������������       �               ��/����?)       *                 �0i?��H\i1�?        �?���J@������������������������       �               ��/����?+       4                 1[v?�x�<�?       �9���*J@,       3                 @*tC?Д�1�B�?       [����D@-       2                 ��c�?P�$3�i�?       ��7���C@.       /                 (�+0?�N:�*ط?       I�G�3@������������������������       �        	       ��,���1@0       1                  <�|?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �        
       ������3@������������������������       �      �<       ��/����?5       8                 �zc?dn����?       � ��w<(@6       7                 pTF�?f%@�"�?       ��[�@������������������������       �               ��#�� @������������������������       �      ��       ��/���@������������������������       �               z�5��@:       I                 pl�{?�]a\��?2       Ut-��xR@;       @                  ��r?k�e���?       �	~�a5@<       ?                    �?4=�%�?       �(J��@=       >                  �P��?bn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               ��/����?A       H                 ���?\O���?       ��o0@B       G                  �JV�?����VV�?
       A�R.�.@C       D                    �?���mf�?       毠�?b@������������������������       �               �cp>@E       F                 H�{�?~�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               鰑%@������������������������       �      �<       ��#���?J       ]                 `���?6x����?"       	V�X@J@K       X                 h���?*4rS7��?       �m��v;@L       Q                 p�s�?�&�+�?	       q��wy�+@M       P                 ��R�?Ȕfm���?       ��Z�N@N       O                 @"@�?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               ��/���@R       S                 0��?�djH�E�?       ^�\m�n@������������������������       �               ��#�� @T       U                 ���?r�T���?       ��e[�&@������������������������       �               ��#�� @V       W                 ��Q�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?Y       \                 �4��?M�#O���?	       �wtJ*@Z       [                 �"��?�_�A�?       炵�e`@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?������������������������       �               H�4H�4@^       g                 �^<:?�T`�[k�?       n��F:l9@_       b                 P�?��Ӭ%�?
       ܅��p3@`       a                  @(B�?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?c       d                    �?�C=+��?       b��T|0@������������������������       �               ��#�� @e       f                 �۲?��=�Sο?       ����,@������������������������       �               ��b:��*@������������������������       �      ȼ       ��/����?h       k                 0v=�?���/��?       @z$S��@i       j                  7u�?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@������������������������       �      м       ��/����?m       n                 `���?�3`���?       .�r��0@������������������������       �               z�5��@o       v                 0/h�?֘�?ʊ�?       ��l���)@p       q                 pʻ�?���3�?       &��X&@������������������������       �               ��+��+@r       s                    �?������?       ���'��@������������������������       �               H�4H�4@t       u                  P���?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ȼ       ��/����?x       �                 p�:?��P�>�?       ԍ�R%(@@y       ~                 ���?* k�Lj�?       e*�}#<=@z       {                 �M�|?^�T��?       ��R�)@������������������������       �               0����/@|       }                 �j%�?<9�)\e�?       _���b @������������������������       �               �cp>@������������������������       �               ;��,��@       �                 `7h�?x�i�@M�?       ���wzb0@������������������������       �               ��/���.@������������������������       �      �<       ��#���?�       �                 ;��?H����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @�       �                 :�?(��_��?       ��B��eH@�       �                 `��?��=��>�?       �n#?4A@�       �                 P2�?�.:�c�?       �Ol2 :@�       �                 p��?\�E�,�?       �MI9@�       �                 �b��?�����o�?       ]���v<3@������������������������       �        
       E�JԮD1@�       �                 �z;y?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                    �?��íxq�?       $2��-�@�       �                  �{?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@�       �                 �7�?v�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0#�?�       �                 GҎi?      �<       ��#�� @������������������������       �               ��#��@������������������������       �               ��#��@�       �                 PT��?      �<	       ��|��,@������������������������       �               ��/����?������������������������       �               ��On�(@�       �                 �}�?��.G��?"       ���\ H@�       �                    �?wT �+��?       ��>Y��@�       �                 �r�?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               �cp>@�       �                 p�?���ճC�?       鰑E@�       �                 h~��?`�ih�<�?       W�3D*5@�       �                 0�!�?8L�0�h�?       l�e�3@������������������������       �               H�4H�4(@�       �                 �+�[?d�ih�<�?       ��
@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                 �n�?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?�       �                 �$I�?      �<       ��-��-5@������������������������       �               0#0# @������������������������       �               ��)��)3@�       �                 �'Q�?�+e�`�?Q       ;��+��]@�       �                 ��9}?�(�q�?       S65�B@�       �                 `��?Hd�9��?       {���(x9@�       �                 r���?�iE���?        ��_�8"@�       �                 ����?��V���?       �0��M @�       �                �E9�?|��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �      ��       ;��,��@������������������������       �      ȼ       ��/����?�       �                  MѴ?�)L垽?       |��[0@�       �                  �P��?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �        	       ���-��*@�       �                  �JV�?      �<       H�4H�4(@������������������������       �               0#0# @������������������������       �               ��+��+$@�       �                 �/��?���Oi��?7       �(}��T@�       �                 0MP�?������?+       sț��P@�       �                 p���?�m(b���?       >O���E@�       �                 p�z�?f���~�?       �v����@@������������������������       �               ��+��+$@�       �                 ���?��)n�?       ����7@������������������������       �               �cp>@�       �                 @��?P��
O&�?       ��(	5@�       �                 �	I�?�W�i6�?       �1�~e1@�       �                  �0��?x�]�uJ�?
       ���:O.@������������������������       �               vb'vb'"@�       �                 (�k�?�D�-,�?       �D'ŰO@�       �                 �;�?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               0#0#@�       �                 pl8�?��G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 �*�?Ҕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@�       �                    �?      �<       vb'vb'"@������������������������       �               0#0# @������������������������       �               �C=�C=@������������������������       �               H�4H�48@�       �                 ��{�?ȇ��?       ��8.@������������������������       �               ��#���?�       �                 P:{�?���!��?       �@��&,@�       �                  =�a?;�N9���?	       ��{j�$@�       �                    �?�g�vw�?       �Aws}8@������������������������       �               ��/����?�       �                 ���?    ��?       "F�b@������������������������       �               ��#���?�       �                 �ie�?b,���O�?       ���/>@������������������������       �               H�4H�4@������������������������       �               ��#���?�       �                  ���?����|e�?       �z �B�@�       �                 �n��?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0# @������������������������       �               0#0#@�t�bh�hhK ��h��R�(KK�KK��h �B  cCy��d@d
���c@yb'vb'b@������c@����/�`@.��+��N@��b:��c@^�_���_@��+��+4@��Gp_b@F��t��V@S2%S2%1@k1��tVa@��t�HQ@0#0#0@#�}��`@��P@0#0# @��#��0@%jW�v%4@        ��#��@                {�5��(@%jW�v%4@        z�5��@                z�5��@&jW�v%4@        ��#���?On��O0@        ��#���?�cp>@                �cp>@        ��#���?                        ���-��*@                ��/����?                ��On�(@        ;��,��@��/���@        ;��,��@��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#��@                        �cp>@            �]@h
��F@0#0# @�k(��B@0����/@        �k(��B@�cp>@        ��#��@@��/����?        ��#��@@                        ��/����?        ��#��@��/����?                ��/����?        ��#��@                        ��/����?                ��/����?                ��/����?        ��k(/T@������C@0#0# @����JG@��/���@                ��/����?        ����JG@���-��@                ��/����?        ����JG@�cp>@        e:��,&C@��/����?        e:��,&C@��/����?        �k(��2@��/����?        ��,���1@                ��#���?��/����?        ��#���?                        ��/����?        ������3@                        ��/����?        ��#�� @��/���@        ��#�� @��/���@        ��#�� @                        ��/���@        z�5��@                Ey�5A@�]�ڕ�?@0#0# @z�5��@D�JԮD1@0#0#�?��#�� @�cp>@        ��#�� @��/����?                ��/����?        ��#�� @                        ��/����?        ��#���?��|��,@0#0#�?        ��|��,@0#0#�?        ��/���@0#0#�?        �cp>@                ��/����?0#0#�?        ��/����?                        0#0#�?        鰑%@        ��#���?                �P^Cy?@��|��,@�C=�C=@[Lg1��&@D�JԮD!@�C=�C=@z�5��@���-��@0#0#�?��#�� @�cp>@        ��#�� @��/����?                ��/����?        ��#�� @                        ��/���@        ��#��@��/����?0#0#�?��#�� @                ��#�� @��/����?0#0#�?��#�� @                        ��/����?0#0#�?        ��/����?                        0#0#�?;��,��@��/����?H�4H�4@;��,��@��/����?        ;��,��@                        ��/����?                        H�4H�4@������3@�cp>@        ��#��0@�cp>@        ��#���?��/����?        ��#���?                        ��/����?        �P^Cy/@��/����?        ��#�� @                ��b:��*@��/����?        ��b:��*@                        ��/����?        z�5��@�cp>@        z�5��@��/����?                ��/����?        z�5��@                        ��/����?        ��#��@��/���@0#0# @z�5��@                ��#���?��/���@0#0# @��#���?��/����?0#0# @                ��+��+@��#���?��/����?H�4H�4@                H�4H�4@��#���?��/����?        ��#���?                        ��/����?                ��/����?        ��#�� @�cp>7@0#0#�?z�5��@�cp>7@        ;��,��@��/���@                0����/@        ;��,��@�cp>@                �cp>@        ;��,��@                ��#���?��/���.@                ��/���.@        ��#���?                ��#�� @        0#0#�?                0#0#�?��#�� @                �k(��"@:l��F:B@H�4H�4@�k(��"@h
��6@H�4H�4@��#���?h
��6@H�4H�4@��#���?h
��6@0#0# @        :l��F:2@0#0#�?        E�JԮD1@                ��/����?0#0#�?                0#0#�?        ��/����?        ��#���?��/���@0#0#�?��#���?�cp>@        ��#���?                        �cp>@                ��/����?0#0#�?                0#0#�?        ��/����?                        0#0#�?��#�� @                ��#��@                ��#��@                        ��|��,@                ��/����?                ��On�(@        ��#���?�cp>@�ڬ�ڬD@��#���?�cp>@0#0# @��#���?        0#0# @��#���?                                0#0# @        �cp>@                �cp>@������C@        �cp>@vb'vb'2@        ��/����?vb'vb'2@                H�4H�4(@        ��/����?H�4H�4@        ��/����?                        H�4H�4@        ��/����?                ��/����?                ��/����?                        ��-��-5@                0#0# @                ��)��)3@<��,��$@�cp>�9@�fm�f�T@;��,��@D�JԮD1@�A�A.@;��,��@D�JԮD1@H�4H�4@;��,��@��/����?0#0# @;��,��@��/����?0#0# @        ��/����?0#0# @                0#0# @        ��/����?        ;��,��@                        ��/����?                ��/���.@0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                ���-��*@                        H�4H�4(@                0#0# @                ��+��+$@;��,��@E�JԮD!@V2%S2%Q@��#�� @���-��@�s?�s?M@��#�� @���-��@S2%S2%A@��#�� @���-��@k�6k�69@                ��+��+$@��#�� @���-��@�A�A.@        �cp>@        ��#�� @��/���@�A�A.@��#���?��/����?�A�A.@��#���?        �C=�C=,@                vb'vb'"@��#���?        ��+��+@��#���?        0#0#�?                0#0#�?��#���?                                0#0#@        ��/����?0#0#�?                0#0#�?        ��/����?        ��#���?�cp>@        ��#���?                        �cp>@                        vb'vb'"@                0#0# @                �C=�C=@                H�4H�48@z�5��@��/����?��+��+$@��#���?                ��#�� @��/����?��+��+$@��#�� @��/����?H�4H�4@��#�� @��/����?H�4H�4@        ��/����?        ��#�� @        H�4H�4@��#���?                ��#���?        H�4H�4@                H�4H�4@��#���?                        ��/����?H�4H�4@        ��/����?0#0#�?                0#0#�?        ��/����?                        0#0# @                0#0#@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJg�$hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKh��BH4         �                 p��?�q�M�N�?'      ��F1Ȋ}@                        �`>R?R�BI$p�?�       �7{<�q@                         @�a�?�`@s'��?       Ei_y,*;@                        �]t?)���?       �� �0!:@                        ��IL?44|���?       	�T|qt2@                         P��?j��H��?       v�I�@       
                  @?��?d%@�"�?       ��[�@       	                 0��>`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               �cp>@������������������������       �               ��#���?                        N��S?      �<       �cp>'@������������������������       �               E�JԮD!@������������������������       �               �cp>@������������������������       �               ��/���@������������������������       �      �<       ��#���?       [                    �?
枞N	�?�       c$���p@       Z                 0!�e?^y,�:��?^       ���ڧyc@       S                 ��z?F����?Y       i3���b@                         �^��?n��H���?I       �,�!�H_@                        8���?jQ��?       �s�=�!@                        P��F?h�r{��?       e�6� @                         `Lվf%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �               0����/@������������������������       �               ��#���?       P                  �m?� �J���?B       3~e]@       3                 P�hf?�\FW��?>       ���Z@       $                 `("?�(߫$��?#        M@~�P@        !                 0��>p)��ĭ?       ��[��@@������������������������       �               ��#��0@"       #                 ��h�>(k� ѽ?	       �����.@������������������������       �               ��/����?������������������������       �               ���>��,@%       0                 �a�?��w���?       W�$�sAA@&       /                 �/��?�����?       �h�d��>@'       ,                 �ЌT?�M:���?
       ����71@(       +                   ��?�����?       �O��(@)       *                 �?����X��?       &��֞&@������������������������       �      ��       ;��,��$@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?-       .                 �+>\?4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @������������������������       �               ��b:��*@1       2                  PV��?      �<       ��/���@������������������������       �               ��/����?������������������������       �               �cp>@4       5                 �T�g?5��`��?       7���?�D@������������������������       �               0#0# @6       A                 `�ռ?"ߩl8�?       U�f�C@7       >                 ��|�?��M��,�?       x��r�0@8       9                 P��?�+�z���?	       LGh��
)@������������������������       �               ��/���@:       ;                  �*x?���mf�?       毠�?b@������������������������       �               ��/����?<       =                   �x�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����??       @                 ����?�zœ���?       IG���t@������������������������       �               0#0#�?������������������������       �               z�5��@B       G                 ��v�?��~'t,�?       ��Ȭc6@C       D                  ���?l7Y���?       ���r�&@������������������������       �               z�5��@E       F                 �/��?L� P?)�?       ����x�@������������������������       �               ��#��@������������������������       �               0#0#�?H       I                  ��?<b����?       �}IS&@������������������������       �               ��#��@J       O                  �6��?n��w��?       ���@K       L                 �j%?��`i��?       �؛.�@������������������������       �               0#0# @M       N                  ���?f%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �      �<       ��/����?Q       R                 𩞺?vQ��?       �s�=�!@������������������������       �               ��#�� @������������������������       �               ���-��@T       U                 �]��?��6L�n�?       ��4}i�8@������������������������       �               <��,��$@V       W                 �u?�B���?       F��,�,@������������������������       �               ��/����?X       Y                 @�:�?lb8�Y�?	       FJͰ(@������������������������       �               ��/����?������������������������       �      �<       [Lg1��&@������������������������       �     �
�       H�4H�4@\       �                  \?�'��u0�??       ��Y@]       f                   ҏ�?j���O�?2       �IR9xKR@^       a                  
?�L����?       [k���>)@_       `                  �Ԧ�?      �<       ��/���@������������������������       �               ��/����?������������������������       �               �cp>@b       e                 �5W�?
4=�%�?       �(J��@c       d                 ��=�?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      �<       ��/����?g       �                 �2OF?v�U���?+       �x�K1GN@h       {                 �$�?����?%       �L�k�nI@i       z                 �{��?�������?       ��4 ��C@j       s                 н��?bn����?       � ��w<8@k       p                 @F�LF�X��?       -�=k�U0@l       o                 @�>\n����?       � ��w<@m       n                  ��^�?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               ��#�� @q       r                 0I��?�FO���?       �ߌ$@������������������������       �               �k(��"@������������������������       �      ȼ       ��/����?t       y                  `s�?Jǵ3���?       �q�ͨ�@u       v                 �-�?��|��?       ���ĺw@������������������������       �               ��#���?w       x                 ��ҥ?t@ȱ��?       om���S@������������������������       �               0����/@������������������������       �               ��#���?������������������������       �               ��#���?������������������������       �               �P^Cy/@|       }                 ���?xY�]���?       ��r-4&@������������������������       �               H�4H�4@~       �                  s��?r�T���?       ��e[�& @       �                 Ly�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 ����?�djH�E�?       ^�\m�n@������������������������       �               ��/����?�       �                 `���?L� P?)�?       ����x�@������������������������       �               ��#�� @�       �                  �c�?T����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @�       �                  �u��?���mf�?       寠�?b#@������������������������       �               ��/���@������������������������       �               0#0# @�       �                  �~��? �)�n�?       �b�}{.;@�       �                 �ON�?X�ih�<�?       ��
@������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?������������������������       �        	       ��+��+4@�       �                 ���?W�
����?w       �l�g@�       �                  4�?���z��?7       A�/�vT@�       �                   ��?ƶ5�3B�?       "é�b80@�       �                 �5�?��h��?       S�D'�@�       �                 `0��?��ڰ�x�?       �K�f�@�       �                  $��?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               ��#��@������������������������       �               0#0#�?�       �                 P���?d*�'=P�?        �2"@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 �6Sz?���뚸�?,       w>c�hP@�       �                 `�^}?ƻ�ݭ�?"       |lNٯGI@������������������������       �               H�4H�4@�       �                 ���T?�M�|%)�?        I$ˤg�G@�       �                 ���?K��*�?       ��X@A@�       �                   +Y�?^�2����?       7#�F�@@�       �                 ��ǻ?��2uj�?       m溕;@�       �                 ��=�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 `A��?dh�iZ�?       TY���$9@�       �                 ��%�?��Ik���?       ��c��.-@�       �                 �[��?��2uj�?
       l溕+@�       �                 ����?�+�z���?	       LGh��
)@�       �                 �?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �               E�JԮD!@������������������������       �      �<       ��#���?������������������������       �      �<       ��#���?������������������������       �               鰑%@�       �                 ��k�?4=�%�?       �(J��@�       �                 �S�?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               ��#���?�       �                    �?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?�       �                 p��U?      �<       ���-��*@������������������������       �               ��/����?������������������������       �               ��On�(@�       �                 P!d�?P��(v��?
       �A�s(.@������������������������       �               ��8��8*@�       �                 ��?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 �|_�?|w+��?@       ���/�Z@�       �                  ���?|�?]b�?)       ��%��Q@�       �                 �+�[?恸�V/�?
       ����|
*@�       �                 ��0�?
4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @�       �                 �ڡS?����?       �a�E�$ @�       �                 𡔜?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               ��+��+@�       �                  �9��?�SA�8�?       ��Ց�L@������������������������       �               ��#�� @�       �                 �x�?���K�?       xVS��K@�       �                 �؈�?h�Ln���?       ���c��J@�       �                  @���?xdhf��?       /l]�
C@�       �                 ��F�?��Eڷ�?       6�L��B@�       �                  `���?(,N=� �?       ��a��+1@�       �                    �?�D#���?       �B�j@������������������������       �               0#0#�?�       �                 ���?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               �C=�C=,@�       �                 0x6�?*^�yU�?       ��7�1�3@�       �                  ���?�� ��?       rp� k@������������������������       �               0#0#�?�       �                  �8�?���mf�?       毠�?b@������������������������       �      �<       ��/���@������������������������       �               0#0#�?�       �                 @Č�?P�ih�<�?       ��
,@�       �                  k&�?�n���k�?       3��&�*@������������������������       �               ��/����?������������������������       �               H�4H�4(@������������������������       �      ȼ       ��/����?������������������������       �      �<       ��#���?�       �                 �@�?      �<       �A�A.@������������������������       �               H�4H�4@������������������������       �               H�4H�4(@������������������������       �      �<       ��/����?�       �                 �|c�?��D4���?       �!�m.�B@������������������������       �               =�C=�C?@�       �                 p4N�?,y��]0�?       ���y"@������������������������       �               ��/����?������������������������       �               ��+��+@�t�bh�hhK ��h��R�(KK�KK��h �Bh  	��GPd@����Xb@�N��Nld@�}��a@�F:l�CW@&S2%S2G@��#��@�cp>7@        z�5��@�cp>7@        z�5��@��/���.@        z�5��@��/���@        ��#�� @��/���@        ��#�� @��/����?                ��/����?        ��#�� @                        �cp>@        ��#���?                        �cp>'@                E�JԮD!@                �cp>@                ��/���@        ��#���?                |�5�wa@M!��Q@&S2%S2G@�}�\Y@�)�B�D@��8��8*@�}�\Y@�)�B�D@�C=�C=@�b:���S@0����/C@�C=�C=@��#�� @���-��@        ��#���?���-��@        ��#���?��/����?                ��/����?        ��#���?                        0����/@        ��#���?                ���khS@�]�ڕ�?@�C=�C=@B����R@��On�8@�C=�C=@t�}wL@0����/#@        �P^Cy?@��/����?        ��#��0@                ���>��,@��/����?                ��/����?        ���>��,@                �#���9@D�JԮD!@        
�#���9@0����/@        z�5��(@0����/@        ;��,��$@��/����?        <��,��$@��/����?        ;��,��$@                        ��/����?                ��/����?        ��#�� @�cp>@                �cp>@        ��#�� @                ��b:��*@                        ��/���@                ��/����?                �cp>@        �k(��2@��/���.@�C=�C=@                0#0# @�k(��2@��/���.@��+��+@z�5��@�cp>'@0#0# @        �cp>'@0#0#�?        ��/���@                ��/���@0#0#�?        ��/����?                ��/����?0#0#�?                0#0#�?        ��/����?        z�5��@        0#0#�?                0#0#�?z�5��@                �P^Cy/@��/���@H�4H�4@<��,��$@        0#0#�?z�5��@                ��#��@        0#0#�?��#��@                                0#0#�?;��,��@��/���@0#0# @��#��@                ��#���?��/���@0#0# @��#���?��/����?0#0# @                0#0# @��#���?��/����?                ��/����?        ��#���?                        ��/����?        ��#�� @���-��@        ��#�� @                        ���-��@        �k(���5@�cp>@        <��,��$@                \Lg1��&@�cp>@                ��/����?        ZLg1��&@��/����?                ��/����?        [Lg1��&@                                H�4H�4@f:��,&C@��|��<@B�A�@@f:��,&C@�a#6�;@�C=�C=@��#�� @鰑%@                ��/���@                ��/����?                �cp>@        ��#�� @�cp>@        ��#�� @��/����?                ��/����?        ��#�� @                        ��/����?        �YLg1B@D�JԮD1@�C=�C=@�YLg1B@/����/#@��+��+@���b:@@��/���@        ��#��0@��/���@        ��b:��*@�cp>@        ��#��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ��#�� @                �k(��"@��/����?        �k(��"@                        ��/����?        z�5��@0����/@        ��#�� @0����/@        ��#���?                ��#���?0����/@                0����/@        ��#���?                ��#���?                �P^Cy/@                ��#��@��/����?��+��+@                H�4H�4@��#��@��/����?0#0# @        ��/����?0#0#�?        ��/����?                        0#0#�?��#��@��/����?0#0#�?        ��/����?        ��#��@        0#0#�?��#�� @                ��#�� @        0#0#�?                0#0#�?��#�� @                        ��/���@0#0# @        ��/���@                        0#0# @        ��/����?��8��8:@        ��/����?H�4H�4@                H�4H�4@        ��/����?                        ��+��+4@�k(��2@���-��J@�s?�s?]@<��,��$@�)�B�D@�A�A>@;��,��@��/����?��+��+$@;��,��@        0#0# @;��,��@        0#0#�?��#���?        0#0#�?                0#0#�?��#���?                ��#��@                                0#0#�?        ��/����?0#0# @        ��/����?                        0#0# @;��,��@&jW�v%D@��+��+4@;��,��@������C@H�4H�4@                H�4H�4@;��,��@������C@H�4H�4@;��,��@�cp>�9@H�4H�4@��#��@�cp>�9@0#0# @��#�� @�cp>7@0#0# @        ��/����?0#0#�?        ��/����?                        0#0#�?��#�� @h
��6@0#0#�?��#�� @�cp>'@0#0#�?��#���?�cp>'@0#0#�?        �cp>'@0#0#�?        �cp>@0#0#�?        �cp>@                        0#0#�?        E�JԮD!@        ��#���?                ��#���?                        鰑%@        ��#�� @�cp>@        ��#���?�cp>@        ��#���?                        �cp>@        ��#���?                ��#���?        0#0#�?��#���?                                0#0#�?        ���-��*@                ��/����?                ��On�(@                ��/����?�C=�C=,@                ��8��8*@        ��/����?0#0#�?        ��/����?                        0#0#�?��#�� @��On�(@�
��
�U@��#�� @�cp>'@l�6k�6I@��#��@��/���@��+��+@��#�� @�cp>@                �cp>@        ��#�� @                ��#�� @��/����?��+��+@��#�� @��/����?                ��/����?        ��#�� @                                ��+��+@��#��@��/���@;�;�F@��#�� @                ��#�� @��/���@;�;�F@��#�� @�cp>@;�;�F@��#�� @�cp>@�A�A>@��#���?�cp>@�A�A>@��#���?        0#0#0@��#���?        0#0# @                0#0#�?��#���?        0#0#�?��#���?                                0#0#�?                �C=�C=,@        �cp>@�C=�C=,@        ��/���@0#0# @                0#0#�?        ��/���@0#0#�?        ��/���@                        0#0#�?        ��/����?H�4H�4(@        ��/����?H�4H�4(@        ��/����?                        H�4H�4(@        ��/����?        ��#���?                                �A�A.@                H�4H�4@                H�4H�4(@        ��/����?                ��/����?vb'vb'B@                =�C=�C?@        ��/����?��+��+@        ��/����?                        ��+��+@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�>D5hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK߅�h��B�0         �                 pY7e?�T�\MO�?&      ����D�}@       �                 `��?��.Q��?�       嗭̟uv@       �                 p웟?����[��?�       �s�D�%v@       i                 P^N<?��t���?�       pb!:p@       &                 ��l?*vϠ��?y       ߠT�Sh@       	                 0��>RfG��?       ��/�.�I@                        ����>h�r{��?       e�6� @������������������������       �               ��#���?������������������������       �               ���-��@
       !                 ~`��8�,��y�?       ��VF@                           �?�J���?       ��o�go@@                        P�# ?@9�)\e�?       ^���b0@������������������������       �               ��/����?                        `Fe�?�_�A�?
       炵�e`,@                         ���?�����?       �O��(@                       @N��?f%@�"�?       ��[�@������������������������       �               ��/����?                        ܿ�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       �k(��"@������������������������       �      м       ��/����?                          ��?��߭Q��?
       �QVl�0@                        k�?���/��?       @z$S��'@                       ��$Ka?Ȕfm���?       ��Z�N@                         ��g�?���/��?       V��7�@������������������������       �               ��#���?                        h�K?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��/���@������������������������       �               ��#��@������������������������       �      ��       0����/@"       %                  �x��?����X��?       &��֞&@#       $                 �M"@?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �               z�5��@'       H                 p���?�s�V���?Z       6��P�a@(       ;                 ���d?��@5��?&       ���N@)       2                    �?؍-�8I�?       ��X5��D@*       1                 ,*���$G�F	�?       ��J�?@+       .                 �vu�?�����?	       �Ä�>c(@,       -                 0�?      �<       ;��,��@������������������������       �               ��#���?������������������������       �               ��#��@/       0                  �P�?�)z� ��?       �\�@������������������������       �               ��#��@������������������������       �               �cp>@������������������������       �      ��       ������3@3       6                  P���?rP�D�?       �A��P?$@4       5                 �>�?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ;��,��@7       :                 �ޗ?Ĕfm���?       ��Z�N@8       9               ��d��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��/����?<       G                 `U�?�x:o��?       s��L- 4@=       D                    �?rdhf��?
       ~/l]�
3@>       ?                 �j��?ʢ��'�?       �^��$@������������������������       �               ��/����?@       C                 ����?a�ox��?       
c��0 @A       B                 �-�?      �<       �C=�C=@������������������������       �               0#0#�?������������������������       �               H�4H�4@������������������������       �               ��#���?E       F                     �?d*�'=P�?        �2"@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      �<       ��/����?I       d                   Y��?�������?4       x��O�+T@J       ]                  ��?��-�2�?0       ��eu�R@K       X                  �?��$�?*       ���*Q@L       M                 0I��?H���'0�?       �C�� TB@������������������������       �               ZLg1��&@N       O                 �G�s?��o�G�?       :�� sE9@������������������������       �               �k(��"@P       W                      ���/��?       U��7�/@Q       V                 ��:�?���Ѯ�?       ��GQ&@R       U                 `�?���/��?       @z$S��@S       T                  zu�?�Z�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@������������������������       �      м       ��/����?������������������������       �      �<       ;��,��@������������������������       �      ȼ       0����/@Y       Z                 `U�?p)��ĭ?       ��[��@@������������������������       �               ���>��<@[       \                 ���?dn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @^       c                  �0��?FH����?       ��ϭ
*@_       `                  �ʇ?��`i��?       �؛.�@������������������������       �               ��#���?a       b                 �6͓?|�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               ��#�� @e       f                 �=��?��`i��?       �؛.�@������������������������       �               ��/����?g       h                  ��3�?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?j       s                  �Q�?D�=n(Y�?&       Hh��AP@k       r                   +Y�?t	˧�d�?       ,A{:=6@l       o                 ���@?��٤ݸ?       ��<5�84@m       n                 ��˘?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?p       q                 ���>      �<	       :l��F:2@������������������������       �               ��/����?������������������������       �               E�JԮD1@������������������������       �               0#0# @t       w                 �u)�>��f;b�?       �/�eE@u       v                 (~?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@x       �                 �T�x?L�?�U�?       my�I�B@y       z                  �x��?@v�"��?       ���d`7@������������������������       �               ���-��*@{       �                 P�~�?��
+���?       \Zz�+�#@|                          �0�?�d�$���?       �T�f@}       ~                �Ʌ#x?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ��#�� @�       �                 `���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                   B�?���mf�?       毠�?b@������������������������       �               ��/���@������������������������       �      �<       0#0#�?�       �                 �5R�?���Ww�?	       v��4]�,@������������������������       �               �k(��"@�       �                 0vb�?��b�}�?       ���\�@�       �                 ��w�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               ��#�� @�       �                 h�4�?�X��-U�?=       F̏ܮW@�       �                 ���?,��| ��?4       ����S@�       �                 �m�?�zA��J�?)       ��
R!�M@�       �                 �m��?�R��b�?       =7��>@�       �                 �-��?�T�"��?	       ��`2�Z+@������������������������       �               �cp>@�       �                �o|?"�Jg@��?       ��G� �%@�       �                  {@�?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?�       �                    �?�֪u�_�?       ��?�8@�       �                 h�B?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       ��/���@�       �                  k�?��i�@M�?       ���wzb0@�       �                 ����?$ k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?������������������������       �      �<	       �cp>'@�       �                 @If�?�@ї�8�?       ���=@�       �                 �i�?,��~d��?
       6E���*@�       �                 �W�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       �cp>'@�       �                 �&m�?f[
�ݢ�?	       F_�Ș0@�       �                 ���?_�:�g�?       �ȁ7B�&@������������������������       �               H�4H�4@�       �                 �ߒ�?��t1u�?       "�te!� @������������������������       �               ��#��@�       �                 X�?�zœ���?       IG���t@������������������������       �               z�5��@������������������������       �               0#0#�?������������������������       �               0����/@�       �                 �==�?�'|5�M�?       ��]�3@������������������������       �               H�4H�4@�       �                 �6��?�&�+�?	       p��wy�+@�       �                 ��N�?����?       ��X�)B @������������������������       �               ��/����?�       �                 ��6�?l����?       P	K��@������������������������       �               ��/����?������������������������       �               z�5��@�       �                 tM�D?�֪u�_�?       ��?�8@�       �                 ੒�?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �               ��/����?�       �                 p��!?      �<	       �A�A.@������������������������       �               ��+��+$@������������������������       �               ��+��+@�       �                 (I��? @����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?�       �                  ���?����X �?F       &���V\@�       �                 @�r�?t�N��?       �XH��)@�       �                    �?r@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@�       �                 �ۢ�?      �<       �C=�C=@������������������������       �               0#0#�?������������������������       �               H�4H�4@�       �                 p�Z�?\(.�??       Q��Y@�       �                    �?�6R�!N�?2       +{�`S@������������������������       �               xb'vb'B@�       �                  �E�?p|�����?       
�/���D@�       �                  `��?��AA#�?       �>�:@�       �                  s��?�~���9�?       �q�Ί#6@�       �                 8c�?�@����?       ���a�@�       �                 �"��?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      ��       0#0# @������������������������       �      ��	       S2%S2%1@�       �                 �	ݡ?��G���?       ��%�|@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �      ��	       �A�A.@�       �                 �1a�?f���;)�?       B��"Z�6@������������������������       �               #0#0&@�       �                 @���? ��ό��?       ���C��'@������������������������       �               0����/@������������������������       �               �C=�C=@�t�bh�hhK ��h��R�(KK�KK��h �B�  ?��,��d@��z��wb@�6k�6�c@-�����d@�]�ڕ�`@����M@-�����d@�-����`@�+��+�K@1�����b@��]�ڕU@%S2%S27@�t�Y,`@
�cp>G@��)��)3@*�����;@�e�_��7@        ��#���?���-��@        ��#���?                        ���-��@        ��b:��:@D�JԮD1@        ��#��0@Nn��O0@        <��,��$@�cp>@                ��/����?        ;��,��$@��/���@        ;��,��$@��/����?        ��#���?��/����?                ��/����?        ��#���?��/����?                ��/����?        ��#���?                �k(��"@                        ��/����?        z�5��@鰑%@        z�5��@�cp>@        ��#�� @�cp>@        ��#�� @��/����?        ��#���?                ��#���?��/����?        ��#���?                        ��/����?                ��/���@        ��#��@                        0����/@        ;��,��$@��/����?        ��#��@��/����?                ��/����?        ��#��@                z�5��@                �}�\Y@h
��6@��)��)3@�k(��B@0����/#@�A�A.@�YLg1B@�cp>@        ���>��<@�cp>@        �k(��"@�cp>@        ;��,��@                ��#���?                ��#��@                ��#��@�cp>@        ��#��@                        �cp>@        ������3@                ���>��@�cp>@        z�5��@                ��#���?                ;��,��@                ��#���?�cp>@        ��#���?��/����?        ��#���?                        ��/����?                ��/����?        ��#���?��/���@�A�A.@��#���?�cp>@�A�A.@��#���?��/����?�C=�C=@        ��/����?        ��#���?        �C=�C=@                �C=�C=@                0#0#�?                H�4H�4@��#���?                        ��/����?0#0# @        ��/����?                        0#0# @        ��/����?        ���b:P@��On�(@0#0#@%�}��O@鰑%@0#0# @Lp�}N@D�JԮD!@        ���>��<@��/���@        ZLg1��&@                ��,���1@��/���@        �k(��"@                ��#�� @��/���@        ��#�� @�cp>@        z�5��@�cp>@        z�5��@��/����?                ��/����?        z�5��@                        ��/����?        ;��,��@                        0����/@        �P^Cy?@��/����?        ���>��<@                ��#�� @��/����?                ��/����?        ��#�� @                z�5��@��/����?0#0# @��#���?��/����?0#0# @��#���?                        ��/����?0#0# @        ��/����?                        0#0# @��#�� @                ��#���?��/����?0#0# @        ��/����?        ��#���?        0#0# @                0#0# @��#���?                <��,��4@'jW�v%D@0#0#@��#���?0����/3@0#0# @��#���?0����/3@        ��#���?��/����?                ��/����?        ��#���?                        :l��F:2@                ��/����?                E�JԮD1@                        0#0# @������3@鰑5@0#0# @��#��@��/����?                ��/����?        ��#��@                �P^Cy/@%jW�v%4@0#0# @��#��@;l��F:2@0#0#�?        ���-��*@        ��#��@0����/@0#0#�?��#��@��/����?        z�5��@                ��#���?                ��#�� @                ��#���?��/����?                ��/����?        ��#���?                        ��/���@0#0#�?        ��/���@                        0#0#�?[Lg1��&@��/����?0#0#�?�k(��"@                ��#�� @��/����?0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?        ��#�� @                ���>��,@�e�_��G@0#0#@@���>��,@�e�_��G@S2%S2%1@��#�� @�)�B�D@��+��+$@��#���?�e�_��7@��+��+@        E�JԮD!@��+��+@        �cp>@                �cp>@��+��+@        ��/����?0#0#@                0#0#@        ��/����?                0����/@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/���@        ��#���?��/���.@        ��#���?��/���@                ��/���@        ��#���?                        �cp>'@        ���>��@E�JԮD1@��+��+@        ��On�(@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>'@        ���>��@0����/@0#0#@���>��@        0#0#@                H�4H�4@���>��@        0#0#�?��#��@                z�5��@        0#0#�?z�5��@                                0#0#�?        0����/@        z�5��@���-��@�C=�C=@                H�4H�4@z�5��@���-��@0#0#�?z�5��@��/����?                ��/����?        z�5��@��/����?                ��/����?        z�5��@                        0����/@0#0#�?        �cp>@0#0#�?        �cp>@                        0#0#�?        ��/����?                        �A�A.@                ��+��+$@                ��+��+@        ��/����?0#0#@                0#0#@        ��/����?        ��#���?��On�(@f'vb'�X@��#���?0����/@�C=�C=@��#���?0����/@        ��#���?                        0����/@                        �C=�C=@                0#0#�?                H�4H�4@        ��/���@,S2%S2W@        �cp>@�z��z�R@                xb'vb'B@        �cp>@��)��)C@        �cp>@%S2%S27@        ��/����?��-��-5@        ��/����?0#0#@        ��/����?0#0# @        ��/����?                        0#0# @                0#0# @                S2%S2%1@        ��/����?0#0# @                0#0# @        ��/����?                        �A�A.@        0����/@vb'vb'2@                #0#0&@        0����/@�C=�C=@        0����/@                        �C=�C=@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ���&hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK˅�h��Bh,         �                 0��v?7]�JU�?/      ��F�\�}@       �                  0C�?�6�$��?�       i7F�fx@       d                 ��~?��c6)T�?�       UmmgO^n@       M                 PUҦ?$S��i/�?y       �/Bl�Xf@                        ��l?�Xm:��?^       5nҟ�/a@                         .:q?��R ��?       +�p�D@                        ���?,µ*A
�?       Su�,h)C@                         Kr6?� �_rK�?       J�@��"@	       
                 ����?�����?       �O��@������������������������       �               ��/����?������������������������       �               ;��,��@������������������������       �               �cp>@                        ��-�?������?        ���O=@������������������������       �               ��#��@                        �o?� ����?       �	��+9@                        H)�[?D3#܅�?       ���A�0@������������������������       �      ��       ��On�(@                        P23? ����?       ��X�)B@                        �p�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?                        .�X?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?                         �0��?      �<       E�JԮD!@������������������������       �               �cp>@������������������������       �               �cp>@                        0H�r?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ��#�� @       @                    �?ڜ����?@       T����X@        5                 �s?fvl6��?.       �:�h�P@!       2                 ��@�?$_蹽�?       �Ǣ�9H@"       1                 @F�h�j���?       �HI�G@#       $                 P��{?�6�x�R�?       ���(�E@������������������������       �        
       ��,���1@%       *                 ��?�d�$���?       	�ٝ9@&       )                 0��_?���/��?       @z$S��@'       (                 �S�?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@������������������������       �      �<       ��/����?+       .                  ��0#����?       x�߄�3@,       -                  `%+�?`n����?       � ��w<@������������������������       �               ��#��@������������������������       �      �<       ��/����?/       0                 p���?      �<
       ��b:��*@������������������������       �               ��#���?������������������������       �        	       z�5��(@������������������������       �               z�5��@3       4                 ��K�?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?6       9                 жd|?���/��?       �[[�.�1@7       8                 p��U?l@ȱ��?       nm���S@������������������������       �      ��       0����/@������������������������       �               ��#���?:       ?                 .w�S?`n����?
       � ��w<(@;       <                 ���@?�d�$���?       �T�f$@������������������������       �      �<       ���>��@=       >                �
�s?Z%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �      м       ��/����?A       F                 P�_!?N��h���?       k��:�=@B       E                   ��?fQ��?       �s�=�!@C       D                 `UMz?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      ��       0����/@G       H                 �2*�?\n����?       ����45@������������������������       �               ��/����?I       L                 �H�=?�����?       ��/̸I3@J       K                 ��N�?k� ѽ?	       �����.@������������������������       �      �<       ���>��,@������������������������       �      ȼ       ��/����?������������������������       �      м       ��/���@N       S                   �P�?�j��?       ��1g�D@O       R                 �=��?�`@s'��?	       Di_y,*+@P       Q                 �}P�?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ȼ       /����/#@T       Y                 `Fe�?�;�F��?       �V�&��;@U       V                 �7ڶ?d*�'=P�?        �2"@������������������������       �               ��+��+@W       X                  �K�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@Z       ]                   �0�?n+}1�?       Vc��2@[       \                 `�"�?�@����?       ���a�@������������������������       �               ��/����?������������������������       �               0#0#@^       c                 ��Q?��n��?       �-H�\+@_       `                    �?�֪u�_�?       ��?�8'@������������������������       �               ��/���@a       b                 X��?z�G���?       ��%�|@������������������������       �      �<       ��/����?������������������������       �               0#0# @������������������������       �               ��#�� @e       |                 �5R�?�-7 
(�?*       n{V�P@f       {                  ��?�Rfv}m�?"       n𼛏I@g       p                 �q*�?&�Rљ�?!       ]�n��I@h       o                 ��ڀ?����ӱ�?       � sE�.0@i       j                 �p�?�B���?       F��,�,@������������������������       �               ���>��@k       l                  �u��?�)z� ��?       �\�@������������������������       �               ��#�� @m       n                 Pm�}?
4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @������������������������       �      м       ��/����?q       z                  S��?����X��?       �f�� �@@r       w                 `Z�?�C=+��?       c��T|@@s       v                 @6�w?\n����?       � ��w<@t       u                 @�:�?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �      ȼ       ��/����?x       y                 �'Yu?      �<       ��b:��:@������������������������       �               ��#�� @������������������������       �               |�5��8@������������������������       �      �<       ��/����?������������������������       �     ��<       0#0#�?}       �                  �_�?�~��v��?       ���*@~                         �a�?��n��?       �-H�\@������������������������       �      ��       0����/@�       �                 ��7�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �      �<       z�5��@�       �                 ��?��E��h�?W       ���mb@�       �                 �p�?*XU�^�?@       "��x�[@�       �                  �~��?�v���?       B��K@@�       �                 `�ܤ?�@G���?	       hu��/@������������������������       �               0#0#@������������������������       �               �cp>'@�       �                 �\�?��i���?       ����1@������������������������       �               ��/����?�       �                 Px��?r����?
       Qz�i0@������������������������       �      ��	       �A�A.@������������������������       �      ȼ       ��/����?�       �                 ��?�?s���?,       稖�S@�       �                 �^Ҧ?_�̣�?%       b�X)P@�       �                  �?b�N�?       �Ȓ���2@�       �                  v_�?����p��?	       �˰�\C+@�       �                 p�3G?�>s{Ab�?       aI��n'@�       �                 ��0�?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �               0����/@������������������������       �               �cp>@�       �                  �-�?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?������������������������       �      �<       ;��,��@�       �                 ��Pw?���o�^�?       �_a�e�F@������������������������       �               H�4H�4@�       �                  h��?(�}���?       �ޗhE@�       �                 `7h�?�~��i9�?       ����\C@�       �                  �u��?P!����?       w��^^A@�       �                 0G�@?x�i�@M�?       ���wzb@@�       �                 ��s'?�3+�Pr�?       [-"�=L4@�       �                 Z&�?� N��?       �L�EBC3@�       �                  �u��?      �<       ���-��*@������������������������       �               ��/����?������������������������       �               �cp>'@�       �                 �1��?l@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@������������������������       �      �<       ��#���?������������������������       �               ��On�(@�       �                  ��?��G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 �3T�?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @�       �                 pH�?�J���?       ��*]Y@������������������������       �               0#0# @������������������������       �               ��#�� @�       �                 p[͔?���i!��?       (��5�,@�       �                 @}�?f,���O�?       ԥ��G](@������������������������       �               0#0# @�       �                  �Ԧ�?�zœ���?       IG���t@������������������������       �               z�5��@������������������������       �               0#0#�?������������������������       �               ��#�� @�       �                  `���?�S�/J�?       ��"Wg�A@�       �                  X3�?�}/W�?       �r�.�%@������������������������       �               ���-��@������������������������       �      ��       0#0#@�       �                 ���?��g�?       ��ʖ�09@������������������������       �               ��/����?�       �                  ���?��E���?       �3q�N;8@�       �                   ���?�k��?       �0QqX@������������������������       �               ��#���?������������������������       �               H�4H�4@������������������������       �        
       S2%S2%1@�       �                 `I9�? �t�Dȗ?5       }"�(iT@�       �                 P�1�?Hy��]0�?       ���y"@������������������������       �               ��+��+@������������������������       �      ȼ       ��/����?������������������������       �      ��/       �i��R@�t�b�     h�hhK ��h��R�(KK�KK��h �B  ��b:��c@�z����c@�6k�6�c@��b:��c@�JԮDmc@������S@Gy�5a@�'�xr�V@0#0#0@�k(���U@�JԮDmS@�C=�C=,@>��,��T@\�v%jWK@        �P^Cy/@�cp>�9@        z�5��(@�cp>�9@        ;��,��@��/���@        ;��,��@��/����?                ��/����?        ;��,��@                        �cp>@        ���>��@h
��6@        ��#��@                z�5��@h
��6@        z�5��@���-��*@                ��On�(@        z�5��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                ��#���?                ��#���?                        E�JԮD!@                �cp>@                �cp>@        z�5��@                ��#���?                ��#�� @                #�}��P@��|��<@        �}�\I@��/���.@        =��,��D@���-��@        >��,��D@0����/@        f:��,&C@0����/@        ��,���1@                <��,��4@0����/@        z�5��@�cp>@        z�5��@��/����?                ��/����?        z�5��@                        ��/����?        ��,���1@��/����?        ��#��@��/����?        ��#��@                        ��/����?        ��b:��*@                ��#���?                z�5��(@                z�5��@                        ��/����?                ��/����?                ��/����?        �k(��"@D�JԮD!@        ��#���?0����/@                0����/@        ��#���?                ��#�� @��/���@        ��#�� @��/����?        ���>��@                ��#���?��/����?                ��/����?        ��#���?                        ��/����?        ��#��0@���-��*@        ��#�� @���-��@        ��#�� @��/����?        ��#�� @                        ��/����?                0����/@        ���>��,@���-��@                ��/����?        ���>��,@0����/@        ���>��,@��/����?        ���>��,@                        ��/����?                ��/���@        ��#��@�cp>7@�C=�C=,@��#�� @�cp>'@        ��#�� @��/����?                ��/����?        ��#�� @                        /����/#@        ��#�� @�cp>'@�C=�C=,@        ��/����?0#0# @                ��+��+@        ��/����?H�4H�4@        ��/����?                        H�4H�4@��#�� @鰑%@H�4H�4@        ��/����?0#0#@        ��/����?                        0#0#@��#�� @0����/#@0#0# @        0����/#@0#0# @        ��/���@                ��/����?0#0# @        ��/����?                        0#0# @��#�� @                ~�5��H@��On�(@0#0# @���#8E@��/���@0#0#�?���#8E@��/���@        ZLg1��&@0����/@        [Lg1��&@�cp>@        ���>��@                ��#��@�cp>@        ��#�� @                ��#�� @�cp>@                �cp>@        ��#�� @                        ��/����?        �P^Cy?@�cp>@        �P^Cy?@��/����?        ��#��@��/����?        ��#��@��/����?                ��/����?        ��#��@                        ��/����?        ��b:��:@                ��#�� @                |�5��8@                        ��/����?                        0#0#�?���>��@0����/@0#0#�?��#���?0����/@0#0#�?        0����/@        ��#���?        0#0#�?��#���?                                0#0#�?z�5��@                ������3@Pn��OP@?�C=�CO@�k(��2@��|��L@fJ�dJ�A@        ���-��*@��)��)3@        �cp>'@0#0#@                0#0#@        �cp>'@                ��/����?�A�A.@        ��/����?                ��/����?�A�A.@                �A�A.@        ��/����?        �k(��2@h
��F@0#0#0@��b:��*@h
��F@�C=�C=@���>��@鰑%@0#0#�?��#�� @鰑%@0#0#�?        鰑%@0#0#�?        0����/@0#0#�?                0#0#�?        0����/@                �cp>@        ��#�� @                ��#���?                ��#���?                ;��,��@                z�5��@�-����@@H�4H�4@                H�4H�4@z�5��@�-����@@H�4H�4@��#��@�-����@@0#0#�?��#�� @�]�ڕ�?@0#0#�?��#�� @��/���>@        ��#�� @;l��F:2@        ��#���?:l��F:2@                ���-��*@                ��/����?                �cp>'@        ��#���?0����/@        ��#���?                        0����/@        ��#���?                        ��On�(@                ��/����?0#0#�?        ��/����?                        0#0#�?��#�� @��/����?                ��/����?        ��#�� @                ��#�� @        0#0# @                0#0# @��#�� @                ;��,��@        vb'vb'"@z�5��@        vb'vb'"@                0#0# @z�5��@        0#0#�?z�5��@                                0#0#�?��#�� @                ��#���?��/���@�;�;;@        ���-��@0#0#@        ���-��@                        0#0#@��#���?��/����?%S2%S27@        ��/����?        ��#���?        %S2%S27@��#���?        H�4H�4@��#���?                                H�4H�4@                S2%S2%1@        ��/����?��+��+T@        ��/����?��+��+@                ��+��+@        ��/����?                        �i��R@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�EhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK���h��B�)         �                 ���? �f$WL�?1      �-P8s}@       �                 `�2|?�D�!��?�       �ՀՕ9w@       p                 p웟?�|v᪣�?�       �N4w&t@       Q                 �� <?�!���s�?�       �P�	p@       N                 �,�?����R�?}       ef�E?7h@       =                 ~`����k���?k       ��X̰c@       8                 H�Y�?9۟qHG�?B       �b�:�W@                        pF�T?]n���2�?>       GX-�[�U@	                        ��`?�^�#΀�?       x�9���?@
                        �J ?xf�T6|�?       z,*��P+@                        �؉�?���/��?       @z$S��@������������������������       �               ��/����?                        �$?Z?����?       ��X�)B@                         h��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?                        �Q�?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?������������������������       �      �<       ��/���@������������������������       �        	       :l��F:2@                        ��j?������?*       V��V�K@������������������������       �        	       <��,��$@                        �~�?�S)D&�?!       ���Km�F@                         �P�?�o���?       o�9�F@                        �xF�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               H�4H�4@       +                  �Q�?|�:�c��?       ��_D��C@       $                 �C8�?��!qP�?       )�9^#�8@        !                 B�F�?jP�D�?       �A��P?$@������������������������       �               ��#��@"       #                 �$I�?���/��?       @z$S��@������������������������       �               �cp>@������������������������       �               z�5��@%       *                 ��Z�?�G��vv�?	       �h� � -@&       '                    �? ��c`�?       &��t5)@������������������������       �               ��/���@(       )                 P�ӕ?* k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?������������������������       �               0#0# @,       5                 �	I�?�K$e_�?       �EU�}.@-       4                 ���r?L[�Jg�?
       X�S0f�*@.       3                 NK�X?��oR��?	       l�Q6�(@/       2                 ��Z�?$�b���?       �GXvƒ@0       1                 �%�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      �<       ;��,��@������������������������       �      ��       ;��,��@������������������������       �      ȼ       ��/����?6       7                 �#��?v�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?9       <                 ��ΐ?0����?       P	K��@:       ;                 ��4�?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               ��#��@>       E                 ��u?@1`f+q�?)       6�W���O@?       @                 p��?�(1k��?       �ꁞ9�F@������������������������       �               ,�����;@A       B                 ue?�x�<�?       X&b��q1@������������������������       �               ��/����?C       D                 O���?�C=+��?       a��T|0@������������������������       �      ��
       �P^Cy/@������������������������       �      ȼ       ��/����?F       I                    �?n%@�"�?
       �6�E�1@G       H                 �j%?      �<       0����/#@������������������������       �               ��/����?������������������������       �               E�JԮD!@J       K                 �5W�?����?       ��X�)B @������������������������       �               z�5��@L       M                ��	��?�Z�	7�?       j~���@������������������������       �               z�5��@������������������������       �      �<       ��/����?O       P                  �{��?0gR���?       ����B@������������������������       �               ��,���A@������������������������       �     ��<       0#0#�?R       m                  �^��?��"m��?,       ܦ�m}pO@S       j                 `���?�`�|���?(       ��6FV\L@T       g                 �2*�?ΫE`P�?#       mT�Ǘ�H@U       \                  �E�?>,���?       �,5��@@V       Y                 �n�]?vf�T6|�?       y,*��P+@W       X                 @F�      �<       0����/#@������������������������       �               ��/���@������������������������       �               ��/����?Z       [                А]�G?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@]       `                 ���?�D���#�?       �C�X��2@^       _                 '4�h?lutee�?       Q9��@������������������������       �               ��/����?������������������������       �               H�4H�4@a       f                 ��>�? :�u���?
       �j7"�5+@b       e                 �6F�?�F���?	       :�.�-'@c       d                  Pmj�?f%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �      ��       D�JԮD!@������������������������       �               0#0# @h       i                 @�V�?�����?
       �N0gX1@������������������������       �      ��	       On��O0@������������������������       �      �<       ��#���?k       l                   ��?�����?       P	K��@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?n       o                �|�?x����1�?       ��;9�@������������������������       �               ��#��@������������������������       �               0#0# @q       �                  ��^�?Ls�DJ��?+       ��dqP@r       y                 ��0�?Dزž �?       ��0(AG@s       x                  ���?�5JH���?       �MOI3@t       u                  y��?H-����?       hM��F2@������������������������       �        
       ��|��,@v       w                 �1��?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �               0#0#�?z       }                  �.�?�(B`P��?       ��A9;@{       |                 @�K?�o���?       o�9�F@������������������������       �               ��#���?������������������������       �               0#0#@~       �                 `}��?F6GzZ��?       �0���'6@       �                 P8��?V�b�z��?       F���2@�       �                 �$��?�@����?       ���a�#@������������������������       �               0#0#@�       �                 �/��?z��`p��?       �����@������������������������       �               ��/����?������������������������       �      ��       0#0#@�       �                 ��?��� ��?       �^�� @������������������������       �               ��/����?�       �                  ��?�djH�E�?       _�\m�n@�       �                  �g<�?      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@�       �                 `<D�?x�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 08��?      �<       ��#��@������������������������       �               ��#�� @������������������������       �               ��#�� @�       �                 ��F�?� N��?       �L�EBC3@������������������������       �               ;l��F:2@������������������������       �      �<       ��#���?�       �                    �?�l
G�f�?        9d�j�H@������������������������       �               H�4H�48@�       �                 P��?�w��Z��?       �R9@������������������������       �        
       �C=�C=,@�       �                 j��?�'z�3�?       ���da�%@������������������������       �               H�4H�4@�       �                 �B��?���mf�?       寠�?b@������������������������       �      ��       ��/���@������������������������       �               0#0#�?�       �                 �dY�?8��ѵ�?>       �_=��X@�       �                 `��?%�C[�?       �;\�9@�       �                 ���?D0�8���?
       #Z��!�)@�       �                 ����?����|e�?	       8\@��'@�       �                  4��?�?�0�!�?       a`�T�$@������������������������       �               ��/����?������������������������       �               vb'vb'"@������������������������       �      ȼ       ��/����?������������������������       �      м       ��/����?�       �                 ����?�����?
       �l�C�J)@�       �                 `��?�n�l���?	       ���5F'@������������������������       �               ��#���?�       �                 �k��?�}	;	�?       vK�>4%@������������������������       �               0����/#@������������������������       �               0#0#�?������������������������       �               0#0#�?�       �                 ���?~��J���?*       g�챂R@�       �                 #s�?f����?       ��F{��J@�       �                  �3��?Hf��{�?       ��C&=@������������������������       �               ��/����?�       �                  P�?����԰?       �����0<@������������������������       �               ��/����?������������������������       �               �;�;;@�       �                 �|'�?lutee�?       �ǟf��8@�       �                 `RZ�?� ����?
       Ӧ����2@������������������������       �               �C=�C=@�       �                  ����?�֪u�_�?       ��?�8'@�       �                    �?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               D�JԮD!@������������������������       �               H�4H�4@�       �                 P�M�?      �<       ��+��+4@������������������������       �               0#0#�?������������������������       �               ��)��)3@�t�bh�hhK ��h��R�(KK�KK��h �B�  C����b@����9e@�����b@1�����b@[<�œb@��)��)S@1�����b@�|�Ǡa@=�C=�C?@}�5�wa@�D�J�.Y@0#0#0@�P^Cy_@;��18N@vb'vb'"@�GpAV@<��18N@0#0# @������C@��h
�G@0#0# @��#��@@�cp>G@0#0# @z�5��@��|��<@        z�5��@鰑%@        z�5��@�cp>@                ��/����?        z�5��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                ��#���?                ��#���?                        ��/���@                :l��F:2@        Lp�}>@E�JԮD1@0#0# @<��,��$@                ������3@D�JԮD1@0#0# @��#���?        0#0#@��#���?        0#0#�?��#���?                                0#0#�?                H�4H�4@�k(��2@D�JԮD1@0#0#@��#�� @��|��,@0#0# @���>��@�cp>@        ��#��@                z�5��@�cp>@                �cp>@        z�5��@                ��#���?�cp>'@0#0# @��#���?�cp>'@                ��/���@        ��#���?��/���@                ��/���@        ��#���?                                0#0# @;��,��$@�cp>@0#0# @<��,��$@��/����?0#0#�?<��,��$@��/����?0#0#�?;��,��@��/����?0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?;��,��@                ;��,��@                        ��/����?                ��/����?0#0#�?                0#0#�?        ��/����?        z�5��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ��#��@                ~�5��H@���-��*@        �k(���E@��/����?        ,�����;@                �P^Cy/@��/����?                ��/����?        �P^Cy/@��/����?        �P^Cy/@                        ��/����?        z�5��@�cp>'@                0����/#@                ��/����?                E�JԮD!@        z�5��@��/����?        z�5��@                z�5��@��/����?        z�5��@                        ��/����?        ��,���A@        0#0#�?��,���A@                                0#0#�?�P^Cy/@)jW�v%D@�C=�C=@\Lg1��&@'jW�v%D@��+��+@;��,��@������C@��+��+@��#��@�cp>7@��+��+@z�5��@鰑%@                0����/#@                ��/���@                ��/����?        z�5��@��/����?                ��/����?        z�5��@                ��#���?��On�(@��+��+@        ��/����?H�4H�4@        ��/����?                        H�4H�4@��#���?鰑%@0#0# @��#���?鰑%@        ��#���?��/����?                ��/����?        ��#���?                        D�JԮD!@                        0#0# @��#���?Pn��O0@                On��O0@        ��#���?                z�5��@��/����?        z�5��@                        ��/����?        ��#��@        0#0# @��#��@                                0#0# @;��,��$@)jW�v%D@�A�A.@�k(��"@h
��6@�A�A.@        D�JԮD1@0#0# @        E�JԮD1@0#0#�?        ��|��,@                �cp>@0#0#�?                0#0#�?        �cp>@                        0#0#�?�k(��"@0����/@��8��8*@��#���?        0#0#@��#���?                                0#0#@��#�� @0����/@vb'vb'"@��#��@0����/@vb'vb'"@        ��/����?0#0# @                0#0#@        ��/����?0#0#@        ��/����?                        0#0#@��#��@�cp>@0#0#�?        ��/����?        ��#��@��/����?0#0#�?��#��@                ��#���?                z�5��@                        ��/����?0#0#�?                0#0#�?        ��/����?        ��#��@                ��#�� @                ��#�� @                ��#���?;l��F:2@                ;l��F:2@        ��#���?                        ��/���@;�;�F@                H�4H�48@        ��/���@��-��-5@                �C=�C=,@        ��/���@�C=�C=@                H�4H�4@        ��/���@0#0#�?        ��/���@                        0#0#�?��#���?��On�8@���~�gR@��#���?���-��*@#0#0&@        ��/���@vb'vb'"@        �cp>@vb'vb'"@        ��/����?vb'vb'"@        ��/����?                        vb'vb'"@        ��/����?                ��/����?        ��#���?0����/#@0#0# @��#���?0����/#@0#0#�?��#���?                        0����/#@0#0#�?        0����/#@                        0#0#�?                0#0#�?        �cp>'@A�C=�CO@        �cp>'@��-��-E@        ��/����?�;�;;@        ��/����?                ��/����?�;�;;@        ��/����?                        �;�;;@        0����/#@�A�A.@        0����/#@vb'vb'"@                �C=�C=@        /����/#@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @        D�JԮD!@                        H�4H�4@                ��+��+4@                0#0#�?                ��)��)3@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ4�phFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKㅔh��B�1         �                  �E�?�+l]>�?(      �����o}@       y                 `�ב?pD4�A��?�       uq��[u@                            �?
��K�?�       ��Y���m@                        ���>�����?       �Һ�b�I@������������������������       �               ��#���?                        p��?�����?       Wb�!�1I@                        �n�?R{��?       �{`g�H@                        ��?��k���?       E+զm7F@	                        �u?r�$�<�?       P���4:@
                        X{e?� ����?       �	��+9@                         ����?* k�Lj�?       d*�}#<-@                        ��?�`@s'��?       Ei_y,*+@������������������������       �               �cp>'@������������������������       �               ��#�� @������������������������       �      �<       ��#���?������������������������       �               鰑%@������������������������       �      �<       ��#���?                        .w�S?      �<	       :l��F:2@������������������������       �               ���-��@������������������������       �               �cp>'@                        ��e�? ���]L�?       N66�ͯ@                        �_��?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �      �<       ��#���?       ^                 �Q��?��#<��?q       4�!+\g@       I                 �+?,����a�?P       ��?�#Q`@       *                 p��a?�Ǩ%���?5       �R �bMV@       %                 @��?��߭Q��?       �QVl�0@       $                 �?9?�_�A�?       肵�e`@        #                 �U�?f%@�"�?       ��[�@!       "                  �P��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      �<       ��/����?������������������������       �               ��#��@&       '                  ��k? ܜ�x�?       d��إV#@������������������������       �               0����/@(       )                  �~��?, k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?+       <                  �_�?�^B��?*       ��k��R@,       7                 pHl?VŠ�T�?       ��0<@-       4                 �!�?�"�Ys��?       ڝ�3@.       3                  Џ~�?�FO���?       �ߌ$@/       0                ���+?�d�$���?       �T�f@������������������������       �      ��       z�5��@1       2                    �?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ;��,��@5       6                   Mt?`Q��?       �s�=�!@������������������������       �               ��#�� @������������������������       �      ��       ���-��@8       ;                 ���R?�"6Aq�?       )$�B"@9       :                 �M��?      �<       �C=�C=@������������������������       �               H�4H�4@������������������������       �               0#0#@������������������������       �      м       ��#�� @=       H                  ��^�?(H�5��?       wqQd� F@>       G                    �?`ڔ>g�?       ���lإE@?       F                 `|\�?�h y/��?       J��.�7@@       A                   s��?����X��?       (��֞6@������������������������       �               ;��,��$@B       C                 P8��?�����?       �O��(@������������������������       �               ���>��@D       E                 �~�?ܗZ�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@������������������������       �               0#0#�?������������������������       �        	       ������3@������������������������       �      �<       ��/����?J       Y                 �Z��?����3#�?       )���ɩD@K       V                  ��d�?��0��~�?       3�3(qA@L       Q                 \F�M?�(���?       �� �0!:@M       N                  ��~�?��/Ѷ?       ���
$6@������������������������       �               ��/���.@O       P                   ��?�`@s'��?       Ei_y,*@������������������������       �               ��#���?������������������������       �               �cp>@R       U                  ����?���/��?       V��7�@S       T                 xb'�?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#���?W       X                 p��Y?F9�)\e�?       _���b @������������������������       �               ;��,��@������������������������       �               �cp>@Z       [                 ��)�?,�b���?       �GXvƒ@������������������������       �               ;��,��@\       ]                 `G,�?x�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?_       p                 P�$�?ȖQ��H�?!       ~m��,L@`       k                 �\��?O�6-�?       lT�ΗD@a       j                  �ف? ꪬD��?       CI)��)>@b       g                 p���?�4�`�?       u�i��]9@c       d                 p�T�?JH����?       ��ϭ
*@������������������������       �               z�5��@e       f                 ���?|�G���?       ��%�|@������������������������       �               0#0# @������������������������       �      �<       ��/����?h       i                  ���?ď%�g�?       ���*wS2@������������������������       �               0#0# @������������������������       �        
       Nn��O0@������������������������       �               0����/@l       m                  �JV�?���3�?       &��X&@������������������������       �               ��#���?n       o                 �c�?�@����?       ���a�#@������������������������       �               ��/����?������������������������       �               0#0# @q       x                 p���?��8��?       Ld\�7Q.@r       w                 0翇?���MF�?       �`�I-*@s       t                 6u�?T������?       "�B(@������������������������       �               vb'vb'"@u       v                 �!�?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �      ȼ       ��/����?������������������������       �               ��#�� @z                         pS��?�#N��F�?C       B���Y@{       |                 pt3�?��t� �?       ����x&@������������������������       �               ��/����?}       ~                 �ڡS?�FO���?       �ߌ$@������������������������       �      ��       �k(��"@������������������������       �      ȼ       ��/����?�       �                 �/Q�?d�)�S[�?=       ��W��W@�       �                 <Ϙ?���D�)�?%       ��@"{wK@�       �                 �)˪?طB" �?       ���<�!*@�       �                  ��d�?|��R[�?       ��"PK&@�       �                 0?�N̸��?       �#�zY9$@������������������������       �               ��#���?������������������������       �               vb'vb'"@������������������������       �      ܼ       ��#���?������������������������       �      ȼ       ��/����?�       �                 �yFC?��h�<*�?       ���D@�       �                  ���?꜋���?       aJ9U63@�       �                 /�?M�����?	       r����.@�       �                 P3"!?      �<       �k(��"@������������������������       �               ���>��@������������������������       �               ��#�� @�       �                 p���?Zn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �      �<       ��/���@�       �                 @�3�?�#:���?       2���ȧ6@������������������������       �               H�4H�4@�       �                  @V��?P+�P���?       �%�8�3@�       �                 ��N�?��^���?       ���w!@�       �                 �Ǒ�?<�a
=�?       ��l��@������������������������       �               0#0#�?������������������������       �               �cp>@�       �                 6u�?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 p���?�'z�3�?
       ���da�%@�       �                  �Ԧ�?|�G���?       ��%�|@������������������������       �               0#0#@������������������������       �      ��       ��/���@������������������������       �               H�4H�4@�       �                   �P�?��/a�N�?       >�n�F�B@�       �                 �D��v=���?       � ��R(@�       �                 p��?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               vb'vb'"@�       �                 �\��?��?'<��?       l��29@�       �                 _%?�s��=��?       ��_��)0@������������������������       �               ��#���?������������������������       �               �A�A.@�       �                 ����?�s:�tp�?       ̾:,"@������������������������       �               ��#��@�       �                 �m��?l�4���?       �tCP��@������������������������       �               �cp>@������������������������       �               0#0# @�       �                 P״�?��eM�?W       3r(`@�       �                   ��?�;�����?       .�3@�       �                 BA�?����|e�?       �z �B�@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?�       �                 P��?ޗZ�	7�?       ���`�$.@�       �                 ��d?���/��?	       ?z$S��'@������������������������       �      ��       z�5��@������������������������       �      ��       �cp>@������������������������       �      ȼ       z�5��@�       �                 @��?����m�?J       �B�V|�[@�       �                 ��ib?x��/���?       ��k�:8?@�       �                 0�!�?��q�R�?       B}Ԥ@������������������������       �               ��/����?�       �                `?��?�J���?       ��*]Y@������������������������       �               ��#�� @������������������������       �               0#0# @������������������������       �      �<       k�6k�69@�       �                 �5Ry?���Aa��?6       &N��m�S@�       �                 ��4�?���S��?$       u��Q�I@�       �                  �P�?��s��/�?       ~��� �B@�       �                  �Mm�?�����?       �O��@������������������������       �               ��#��@�       �                 `�ۊ?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 荤�?����2��?       8���}?@������������������������       �               H�4H�4@�       �                  ���?����N�?       ��G�v<@�       �                 @*��?� ����?       �趩��3@������������������������       �               0����/@�       �                 �Qe�?���(n��?
       b����-@�       �                   ҏ�?D��NV=�?       �t�ܲ@�       �                 P�ͪ?m��w��?       ���@�       �                 @���?�3`���?       .�r��@�       �                   B�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 ��ď?      �<       0#0# @������������������������       �               0#0#�?������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               �C=�C=@�       �                  �u��?<[��G�?	       �O�;�]!@������������������������       �               ��/���@������������������������       �               0#0#�?������������������������       �               �C=�C=,@�       �                 �?�?      �<       �;�;;@������������������������       �               H�4H�4@������������������������       �               H�4H�48@�t�bh�hhK ��h��R�(KK�KK��h �BH  Gy�5a@\�ڕ��d@�fm�f�d@    �]@�|�Ǡa@�ڬ�ڬT@�#����U@A�)�B]@B�A�@@���>��@��]�ڕE@0#0#�?��#���?                z�5��@��]�ڕE@0#0#�?;��,��@��]�ڕE@0#0#�?��#��@&jW�v%D@        ��#��@h
��6@        z�5��@h
��6@        z�5��@�cp>'@        ��#�� @�cp>'@                �cp>'@        ��#�� @                ��#���?                        鰑%@        ��#���?                        :l��F:2@                ���-��@                �cp>'@        ��#���?�cp>@0#0#�?��#���?        0#0#�?                0#0#�?��#���?                        �cp>@        ��#���?                ��k(/T@��z��wR@0#0#@@��Gp_R@�e�_��G@vb'vb'"@Np�}N@鰑5@0#0# @z�5��@鰑%@        ;��,��@��/����?        ��#���?��/����?        ��#���?��/����?        ��#���?                        ��/����?                ��/����?        ��#��@                ��#���?D�JԮD!@                0����/@        ��#���?��/���@                ��/���@        ��#���?                ��b:��J@鰑%@0#0# @��b:��*@��/���@�C=�C=@\Lg1��&@��/���@        �k(��"@��/����?        ��#��@��/����?        z�5��@                ��#���?��/����?        ��#���?                        ��/����?        ;��,��@                ��#�� @���-��@        ��#�� @                        ���-��@        ��#�� @        �C=�C=@                �C=�C=@                H�4H�4@                0#0#@��#�� @                ��k(/D@�cp>@0#0#�?��k(/D@��/����?0#0#�?<��,��4@��/����?0#0#�?<��,��4@��/����?        ;��,��$@                ;��,��$@��/����?        ���>��@                z�5��@��/����?                ��/����?        z�5��@                                0#0#�?������3@                        ��/����?        ��b:��*@���-��:@0#0#�?��#�� @�cp>�9@        z�5��@�cp>7@        ��#���?鰑5@                ��/���.@        ��#���?�cp>@        ��#���?                        �cp>@        ��#�� @��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#���?                ;��,��@�cp>@        ;��,��@                        �cp>@        ;��,��@��/����?0#0#�?;��,��@                        ��/����?0#0#�?                0#0#�?        ��/����?        ���>��@�cp>�9@%S2%S27@��#��@��On�8@H�4H�4(@z�5��@�cp>7@0#0#@z�5��@9l��F:2@0#0#@z�5��@��/����?0#0# @z�5��@                        ��/����?0#0# @                0#0# @        ��/����?                On��O0@0#0# @                0#0# @        Nn��O0@                0����/@        ��#���?��/����?0#0# @��#���?                        ��/����?0#0# @        ��/����?                        0#0# @z�5��@��/����?#0#0&@��#���?��/����?#0#0&@��#���?        #0#0&@                vb'vb'"@��#���?        0#0# @��#���?                                0#0# @        ��/����?        ��#�� @                Jp�}>@�e�_��7@\��Y��H@�k(��"@��/����?                ��/����?        �k(��"@��/����?        �k(��"@                        ��/����?        ;��,��4@h
��6@\��Y��H@�P^Cy/@:l��F:2@��-��-5@��#�� @��/����?vb'vb'"@��#�� @        vb'vb'"@��#���?        vb'vb'"@��#���?                                vb'vb'"@��#���?                        ��/����?        ��b:��*@On��O0@H�4H�4(@��b:��*@�cp>@        ��b:��*@��/����?        �k(��"@                ���>��@                ��#�� @                ��#��@��/����?                ��/����?        ��#��@                        ��/���@                鰑%@H�4H�4(@                H�4H�4@        鰑%@vb'vb'"@        ���-��@0#0# @        �cp>@0#0#�?                0#0#�?        �cp>@                ��/����?0#0#�?        ��/����?                        0#0#�?        ��/���@�C=�C=@        ��/���@0#0#@                0#0#@        ��/���@                        H�4H�4@;��,��@��/���@�C=�C=<@        ��/����?#0#0&@        ��/����?0#0# @        ��/����?                        0#0# @                vb'vb'"@;��,��@�cp>@S2%S2%1@��#���?        �A�A.@��#���?                                �A�A.@��#��@�cp>@0#0# @��#��@                        �cp>@0#0# @        �cp>@                        0#0# @�k(��2@�cp>�9@��-��-U@�k(��"@���-��@H�4H�4@        ��/����?H�4H�4@                H�4H�4@        ��/����?        �k(��"@�cp>@        z�5��@�cp>@        z�5��@                        �cp>@        z�5��@                �k(��"@0����/3@�N��NlT@��#�� @��/����?�;�;;@��#�� @��/����?0#0# @        ��/����?        ��#�� @        0#0# @��#�� @                                0#0# @                k�6k�69@���>��@D�JԮD1@�;�;K@���>��@D�JԮD1@�;�;;@���>��@D�JԮD1@��8��8*@;��,��@��/����?        ��#��@                ��#���?��/����?        ��#���?                        ��/����?        ��#�� @Nn��O0@��8��8*@                H�4H�4@��#�� @On��O0@��+��+$@��#�� @E�JԮD!@vb'vb'"@        0����/@        ��#�� @��/���@vb'vb'"@��#�� @��/���@0#0# @��#���?��/���@0#0# @��#���?��/����?0#0# @��#���?��/����?                ��/����?        ��#���?                                0#0# @                0#0#�?                0#0#�?        �cp>@        ��#���?                                �C=�C=@        ��/���@0#0#�?        ��/���@                        0#0#�?                �C=�C=,@                �;�;;@                H�4H�4@                H�4H�48@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJLxhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKх�h��B�-         �                 pK�b?��)��K�?'      l�⍫�}@       �                 �^Ҧ?ks�:��?�       !{���v@       6                 ��j?�Ҁ�0
�?�       �{�2��q@       3                 P���?2����>�?M       (%�*L]@       *                 �)�?86DU�!�?F       ���^�Z@                         `�J�?4K׀���?A       �#[���X@������������������������       �               ��/����?       )                 �2*�?&�B�y��?@       #d���%X@	                        �U��������'�?5       *RҀh�T@
                        �!}V?��*F��?       j�;=�nA@                        6D�G?h�r{��?       e�6� @������������������������       �               ���-��@������������������������       �               ��#���?                          ��?�$߱�m�?       �}�l?;@                         e	a?|�C<BF�?       ��`��F7@������������������������       �               z�5��@                        �\͵?�\�sF��?       U>��1@                        ����>\����?       P	K��@                        �Q�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ��       ;��,��@                        Ћ�R?
4=�%�?        �(J��#@������������������������       �      ȼ       �cp>@������������������������       �               ��#��@������������������������       �      ��       ��/���@                        ��R?�I��X[�?       �h��G@������������������������       �               ��/����?                        ��L�>\�؈�w�?       q���S#G@������������������������       �               ��/����?       "                 @��>x�+(�s�?       �9Շ�F@        !                  P���?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @#       &                 ��L�?।�N-�?       �#[�$E@$       %                 @*tC?��p?��?       P�^��B@������������������������       �               �YLg1B@������������������������       �      �<       ��/����?'       (                 �IK?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �               ���>��,@+       0                  �?�\z����?       ���U��!@,       -                    �?b,���O�?       ���/>@������������������������       �               0#0# @.       /                 0�!�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?1       2                  ���?& k�Lj�?       �q��l}@������������������������       �               ��/���@������������������������       �      м       ��#���?4       5                  0Y��?��j�Lj�?       �q��l}#@������������������������       �               ��/���@������������������������       �               ��#�� @7       L                 �oz?�|X���?d       ��DP2�d@8       9                 �a ?�]��0�?       ң�Bm�B@������������������������       �               ��#�� @:       I                  `���?ܐ�Q%G�?       Bã�q�A@;       F                 �*U�?�.*���?       �"�t:@<       E                 й�o?@��;��?       �N��b8@=       B                  y��?������?       Wؗյ0@>       ?                 P�\?�F���?	       :�.�-'@������������������������       �               0����/#@@       A                 `��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?C       D                 �\��?�|2N��?       �3K}@������������������������       �               z�5��@������������������������       �               0#0# @������������������������       �               ��/���@G       H                 (�!�?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?J       K                 ȋ�v?      �<       E�JԮD!@������������������������       �               ��/����?������������������������       �               ��/���@M       x                 ���@?PA��9�?K       �;��`@N       k                 `��m?v3,ן��?7       L����W@O       h                 ����?Б�Q���?       ���J@P       [                  @V��?��(�|?�?       Ĝ���wC@Q       X                 �瓠?t����?       ~��qπ*@R       S                 ����?�FO���?       �ߌ$@������������������������       �               ;��,��@T       U                   �G�?~d�$���?       �T�f@������������������������       �               z�5��@V       W                 �{��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?Y       Z                 �U�,?z��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?\       a                  ���?�ѿ�FB�?       H���W�9@]       `                  J��?$ k�Lj�?       �q��l}#@^       _                 �Ix�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ��       ���-��@b       g                 �xȟ?����|e�?	       �z �B�/@c       d                    �?�n���k�?       3��&�*@������������������������       �               vb'vb'"@e       f                  �~��?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �      ȼ       �cp>@i       j                 �vQ?�(߫$��?       1H����*@������������������������       �      �<       [Lg1��&@������������������������       �      ȼ       ��/����?l       w                 �X\�?c��q��?       �Y�r�E@m       v                    �?����?       K�YŦ'E@n       s                  �?�b���:�?
       �
#���,@o       r                 _%?ҟ��X�?       l�n�/@p       q                  h��?�J���?       ��*]Y@������������������������       �               0#0# @������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?t       u                 ���?      �<       �k(��"@������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �               *�����;@������������������������       �      �<       ��/����?y       �                 �=M�?�yoJ	�?       ���8
�@@z       }                 0���?���9��?       ����s4@{       |                �3�r?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @~                        ���?)���?
       y��uk1@������������������������       �      �<       ��On�(@�       �                 �#��?4=�%�?       �(J��@������������������������       �               ��#�� @������������������������       �               �cp>@�       �                 p�O�?������?       y���)@������������������������       �               H�4H�4@�       �                 03�?��|��?       ���ĺw@������������������������       �               ��#���?�       �                    �?r@ȱ��?       om���S@�       �                 �-��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��/���@�       �                  ���?R0��Cb�?0       ��k��hT@�       �                 0�I�?"����?       Ol��PC@�       �                  ��?��&7~��?       ���,A:@�       �                 ��Iz?      �<       0����/3@������������������������       �               ��/����?������������������������       �        
       E�JԮD1@�       �                    �?�26�
�?       5��*8E@�       �                  �g<�?L� P?)�?       ����x�@������������������������       �               z�5��@�       �                 ���?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                  I�?���/��?       ?z$S��'@�       �                 @���?����?       ��X�)B @�       �                 ���?l����?       Q	K��@������������������������       �               ;��,��@�       �                 (�3?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ȼ       ��/����?������������������������       �      м       ��/���@�       �                 ���T?�fa��?       s�7���E@�       �                 0���?�U)m��?       "�$�jdA@�       �                  �.�?��^���?       ���w!@������������������������       �               0#0# @������������������������       �      ��       ���-��@�       �                 0��?x'1n 6�?       E��N:@�       �                 P� �?F�Uέ��?	       Bq��+@������������������������       �               ��/����?�       �                 PeT�?Hj��w�?       l8�(@������������������������       �               H�4H�4@�       �                 ��U�?������?       ���'��@������������������������       �               H�4H�4@�       �                  u��?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �               H�4H�4(@������������������������       �      �       D�JԮD!@�       �                 �=�t?��$�v|�?F       X}��I�Z@������������������������       �               z�5��@�       �                    �?�bJ��i�?E       �T��Z@������������������������       �                ˷|˷I@�       �                   B�?�"��s�?%       X�B�N�J@�       �                 ��O�?�΢~��?       p����C@�       �                 @�ۓ?z�G���?       ��%�|@������������������������       �               ��/���@������������������������       �               0#0#@�       �                 @f�?���L�?       >G���@@������������������������       �               vb'vb'"@�       �                   �?h���;)�?       B��"Z�6@�       �                  ���?�v�;B��?       ՟���	0@�       �                 �3P�?t��ճC�?	       y��l$,@������������������������       �               vb'vb'"@�       �                  ��d�?�@����?       ���a�@������������������������       �               H�4H�4@�       �                 ��?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 @w�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 �81�?�Qk��?       ��Th!�@�       �                 `���?�@G���?       hu��@�       �                 P���?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               H�4H�4@������������������������       �        
       ��8��8*@�t�bh�hhK ��h��R�(KK�KK��h �B�  ���#8e@�JԮDmc@~��~�gb@Qg1���d@����Xb@~˷|˷I@���khc@�D�J�.Y@�;�;;@������S@����z�A@H�4H�4@f:��,&S@�a#6�;@H�4H�4@�k(��R@�e�_��7@                ��/����?        �k(��R@h
��6@        Lp�}N@h
��6@        ��,���1@D�JԮD1@        ��#���?���-��@                ���-��@        ��#���?                ��#��0@鰑%@        ��#��0@���-��@        z�5��@                <��,��$@���-��@        z�5��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ;��,��@                ��#��@�cp>@                �cp>@        ��#��@                        ��/���@        ���#8E@0����/@                ��/����?        ���#8E@��/���@                ��/����?        ���#8E@�cp>@        ��#�� @��/����?                ��/����?        ��#�� @                ��k(/D@��/����?        �YLg1B@��/����?        �YLg1B@                        ��/����?        ��#��@��/����?        ��#��@                        ��/����?        ���>��,@                ��#�� @��/���@H�4H�4@��#���?        H�4H�4@                0#0# @��#���?        0#0#�?��#���?                                0#0#�?��#���?��/���@                ��/���@        ��#���?                ��#�� @��/���@                ��/���@        ��#�� @                f:��,&S@Rn��OP@H�4H�48@��#�� @���-��:@0#0# @��#�� @                z�5��@���-��:@0#0# @z�5��@9l��F:2@0#0# @��#��@9l��F:2@0#0# @��#��@鰑%@0#0# @��#���?鰑%@                0����/#@        ��#���?��/����?                ��/����?        ��#���?                z�5��@        0#0# @z�5��@                                0#0# @        ��/���@        ��#�� @                ��#���?                ��#���?                        E�JԮD!@                ��/����?                ��/���@        Gy�5Q@1����/C@#0#06@�P^CyO@E�JԮD1@0#0#0@[Lg1��6@��/���.@�C=�C=,@\Lg1��&@���-��*@�C=�C=,@�k(��"@��/����?0#0# @�k(��"@��/����?        ;��,��@                ��#��@��/����?        z�5��@                ��#���?��/����?                ��/����?        ��#���?                        ��/����?0#0# @                0#0# @        ��/����?        ��#�� @�cp>'@H�4H�4(@��#�� @��/���@        ��#�� @��/����?                ��/����?        ��#�� @                        ���-��@                ��/���@H�4H�4(@        ��/����?H�4H�4(@                vb'vb'"@        ��/����?H�4H�4@        ��/����?                        H�4H�4@        �cp>@        ZLg1��&@��/����?        [Lg1��&@                        ��/����?        ������C@��/����?0#0# @������C@��/����?0#0# @ZLg1��&@��/����?0#0# @��#�� @��/����?0#0# @��#�� @        0#0# @                0#0# @��#�� @                        ��/����?        �k(��"@                ��#���?                ��#�� @                *�����;@                        ��/����?        z�5��@鰑5@H�4H�4@��#��@On��O0@        ��#�� @��/����?                ��/����?        ��#�� @                ��#�� @��/���.@                ��On�(@        ��#�� @�cp>@        ��#�� @                        �cp>@        ��#�� @0����/@H�4H�4@                H�4H�4@��#�� @0����/@        ��#���?                ��#���?0����/@        ��#���?��/����?        ��#���?                        ��/����?                ��/���@        \Lg1��&@	�cp>G@H�4H�48@;��,��$@���-��:@0#0#�?��#��@鰑5@0#0#�?        0����/3@                ��/����?                E�JԮD1@        ��#��@��/����?0#0#�?��#��@        0#0#�?z�5��@                ��#���?        0#0#�?��#���?                                0#0#�?        ��/����?        z�5��@�cp>@        z�5��@��/����?        z�5��@��/����?        ;��,��@                ��#���?��/����?                ��/����?        ��#���?                        ��/����?                ��/���@        ��#���?0����/3@%S2%S27@��#���?鰑%@%S2%S27@        ���-��@0#0# @                0#0# @        ���-��@        ��#���?��/���@��-��-5@��#���?��/���@vb'vb'"@        ��/����?        ��#���?��/����?vb'vb'"@                H�4H�4@��#���?��/����?H�4H�4@                H�4H�4@��#���?��/����?                ��/����?        ��#���?                                H�4H�4(@        D�JԮD!@        z�5��@D�JԮD!@F�s?��W@z�5��@                        D�JԮD!@B�s?��W@                ˷|˷I@        D�JԮD!@#0#0F@        D�JԮD!@=�C=�C?@        ��/���@0#0#@        ��/���@                        0#0#@        0����/@�;�;;@                vb'vb'"@        0����/@vb'vb'2@        ��/����?�C=�C=,@        ��/����?��8��8*@                vb'vb'"@        ��/����?0#0#@                H�4H�4@        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@0#0#@        �cp>@0#0#�?        �cp>@                ��/����?                ��/����?                        0#0#�?                H�4H�4@                ��8��8*@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJW��8hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKh��BH4         T                 ��{�?C�|���?)      �h���}@       C                 h�l�?��d���?^       k���Eb@       >                 � �l?�����?P       ]7���_@       /                 ��_i?r)�Ug��?F       ��L'��[@                        @�W?�g�Ҥ�?-       	Ǿb4S@       	                  m?��F���?       :�.�-'@                        0��>$ k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?
                        ��L?      �<       ���-��@������������������������       �               ��/����?������������������������       �               0����/@       .                 ߣ�?0Й����?&       �3�NP@                         �P��?�ĕ��F�?%       c7 �S�O@                           �?X ����?
       2
C>�5@������������������������       �               ��b:��*@                        ��_?��6L�n�?       �E#��h @                         ����?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               z�5��@       !                 ��9�?�C$T��?       H����D@                         �M�e?��oR��?       m�Q6�8@                           �?����X��?       (��֞6@                        �F?�#�Ѵ�?       �)�B�4@������������������������       �               ���>��,@                        p��?�����?       �O��@������������������������       �               ��/����?������������������������       �               ;��,��@                        �$I�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               0#0# @"       )                  ��?���Ul��?        {|3�0@#       &                 ���^?lP�D�?       �A��P?$@$       %                 0��>�����?       �O��@������������������������       �               ��/����?������������������������       �               ;��,��@'       (                 �2e?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @*       -                 �Q�?�`@s'��?       Fi_y,*@+       ,                 �U�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               0����/@������������������������       �               0#0# @0       5                  `�J�?�O
�0�?       ���
#A@1       2                    �?�0�~��?       r��GQ1@������������������������       �      ��       ��On�(@3       4                  �"�?���mf�?       寠�?b@������������������������       �      ��       ��/���@������������������������       �               0#0#�?6       7                 l\��?ǋr��?	       ��#���0@������������������������       �               0����/@8       9                 p�p�?Ƴ�F�M�?       S��ڭQ(@������������������������       �               ��#��@:       =                  `���?�v�;B��?       ՟���	 @;       <                  `��?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               H�4H�4@?       B                 @��J?�~�Hs=�?
       ��?Z[0@@       A                  ���?\����?       P	K��,@������������������������       �               z�5��(@������������������������       �      ȼ       ��/����?������������������������       �               0#0# @D       G                 P_RM?�`{���?       �~8�31@E       F                �� ��?�zœ���?       IG���t@������������������������       �               z�5��@������������������������       �               0#0#�?H       S                 ��@�?B0�8���?       "Z��!�)@I       P                 �ߝw?����|e�?       8\@��'@J       K                 `�ܤ?h�4���?       �tCP��@������������������������       �               0#0#�?L       O                 �5��?�@G���?       hu��@M       N                  H��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               0#0#�?Q       R                    �?      �<       �C=�C=@������������������������       �               H�4H�4@������������������������       �               0#0#@������������������������       �      м       ��/����?U       �                 ���?AA!�%.�?�       �rw��t@V       �                 pH�d?8��7c�?Z       eu@^�b@W       z                 �+@?��5O7�?Q       "[��C�`@X       w                 ���?�u��a�?1       lb)~�T@Y       p                 ��N�?�Wߕ�?.       �Q7'T@Z       i                 ��?p^�Y��?       1A���G@[       h                 �V��?�Z�!���?       ��e`��<@\       a                  �ޖ?�Q0TuJ�?       ʃ�Я[5@]       `                 ��kc?��6L�n�?	       �E#��h0@^       _                 ��Z?���/��?       V��7�@������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �      ��       z�5��(@b       e                    �?4=�%�?       �(J��@c       d                 p��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?f       g                   \��?d%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ���>��@j       m                 Aј?r���;��?
       �ڴ���2@k       l                 @C��?$ k�Lj�?       �q��l}#@������������������������       �      ��       ��/���@������������������������       �               ��#�� @n       o                  �\�?H���'0�?       �C�� T"@������������������������       �               ��/����?������������������������       �               ���>��@q       t                 �R�}?�+op�?       ���Ǣr@@r       s                    �?
4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @u       v                    �?      �<       +�����;@������������������������       �               �k(��"@������������������������       �        	       �k(��2@x       y                  �@�?E#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?{       �                   s��?���{�k�?        Y���
J@|       �                   ҏ�?nQ��?       �s�=�1@}       ~                 ��ъ?�)z� ��?       �\�@������������������������       �               ��#�� @       �                    �?
4=�%�?       �(J��@�       �                 ��G�?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      �<       ��/����?�       �                 (]8o?      �<       鰑%@������������������������       �               ��/����?������������������������       �               0����/#@�       �                 ���?����6��?       �Z�K�@A@�       �                 ���?.c{���?       6:���=@�       �                 @')?��6L�n�?       ��4}i�8@������������������������       �               ��/����?�       �                 �H�?���sx�?       �iۍѧ7@�       �                    �?�(1k��?       �ꁞ9�6@������������������������       �               ��#��0@�       �                  ���?�����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?������������������������       �      �<       ��/����?�       �                 ��$j?�������?       "F�b@������������������������       �               ��#�� @������������������������       �               H�4H�4@�       �                 �;ڕ?      �<       0����/@������������������������       �               ��/����?������������������������       �               �cp>@������������������������       �      �	       �A�A.@�       �                   E(�?�(�K��?q       [p��sPf@�       �                 �3ן?:�S-��?       ��-�~�<@�       �                 �T��?�|2N��?       �3K}@������������������������       �               z�5��@������������������������       �               0#0# @�       �                    �?u�%��?       ��l,�7@�       �                 �-�?Ɠ�R �?       ��u�(@������������������������       �               0����/@�       �                 ����? Lj����?       ���T�@�       �                 P�g�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               ;��,��@�       �                 �q
�?      �<	       �cp>'@������������������������       �               ��/����?������������������������       �               鰑%@�       �                 ���?t����?\       �hţ�b@�       �                  �6��?���+1T�?7       �<�8W�V@�       �                 ���?f��oM|�?*       <42�4lQ@�       �                    �?�wƄ(�?       n�V�AG@�       �                 �-�?�Rn*l�?       4���2@�       �                 `��?������?
       ���]�'@������������������������       �               �cp>@�       �                 `�Q�?�\z����?       ���U��!@������������������������       �               ��#���?�       �                  ��?�1�RH3�?       =�����@�       �                 P8��?��íxq�?       %2��-�@������������������������       �               0#0#�?�       �                 �f��?& k�Lj�?       �q��l}@������������������������       �               �cp>@�       �                  `���?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               0#0# @������������������������       �               �C=�C=@�       �                  y�?<���1�?       ��+�N�;@�       �                  ���?�26�
�?       4��*8E,@�       �                 �+3�?l��w��?       ���@�       �                 �_��?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               ��/���@������������������������       �               ���>��@�       �                 �C8�?,e��}�?	       ��Se+@������������������������       �               ��/���@�       �                   �x�?t@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@�       �                 �oo�?z�&�?       �ۄ-7@�       �                  �g<�?L�0�h�?       k�e�3@�       �                 p͹�?�@����?       ���a�@������������������������       �               ��/����?������������������������       �               0#0#@������������������������       �      ��       �C=�C=,@�       �                 �_��?
����?       ��X�)B@������������������������       �               ��#�� @�       �                 �@�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 ��^f?�����?       �!XY�$6@�       �                 �fQ?ַB" �?       ���<�!*@�       �                 pTF�?�o���?       o�9�F$@������������������������       �               ��#�� @������������������������       �               0#0# @�       �                 k�;�?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �               vb'vb'"@�       �                 ����?�Ї�	��?%       LV���M@�       �                 p�?0�-al��?       �h�t}�=@������������������������       �               vb'vb'"@�       �                 ����?FN�\x�?       ���9̶4@�       �                 @��?�;[��G�?       �O�;�]!@�       �                 h��?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �               �cp>@�       �                 p�h�?Rj��w�?       l8�(@�       �                 ���q?��`i��?       �؛.�@�       �                    �?f%@�"�?       ��[�@������������������������       �               ��/����?�       �                  u�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               �C=�C=@������������������������       �      ��       �C=�C=<@�t�b�T     h�hhK ��h��R�(KK�KK��h �Bh  �P^Cy�g@�|�Ǡa@l�fm��a@��,���Q@��On�H@H�4H�48@"�}��P@
�cp>G@�C=�C=,@�>��nK@h
��F@H�4H�4(@�}�\I@h
��6@0#0#@��#���?鰑%@        ��#���?��/���@                ��/���@        ��#���?                        ���-��@                ��/����?                0����/@        |�5��H@�cp>'@0#0#@|�5��H@�cp>'@0#0# @<��,��4@��/����?        ��b:��*@                ���>��@��/����?        ��#���?��/����?                ��/����?        ��#���?                z�5��@                ���>��<@鰑%@0#0# @<��,��4@��/����?0#0# @<��,��4@��/����?        ������3@��/����?        ���>��,@                ;��,��@��/����?                ��/����?        ;��,��@                ��#���?��/����?                ��/����?        ��#���?                                0#0# @��#�� @D�JԮD!@        ���>��@�cp>@        ;��,��@��/����?                ��/����?        ;��,��@                ��#�� @��/����?                ��/����?        ��#�� @                ��#���?�cp>@        ��#���?��/����?                ��/����?        ��#���?                        0����/@                        0#0# @��#��@h
��6@0#0# @        On��O0@0#0#�?        ��On�(@                ��/���@0#0#�?        ��/���@                        0#0#�?��#��@�cp>@�C=�C=@        0����/@        ��#��@��/����?�C=�C=@��#��@                        ��/����?�C=�C=@        ��/����?0#0#�?                0#0#�?        ��/����?                        H�4H�4@z�5��(@��/����?0#0# @z�5��(@��/����?        z�5��(@                        ��/����?                        0#0# @z�5��@��/���@��+��+$@z�5��@        0#0#�?z�5��@                                0#0#�?        ��/���@vb'vb'"@        �cp>@vb'vb'"@        �cp>@0#0# @                0#0#�?        �cp>@0#0#�?        �cp>@                ��/����?                ��/����?                        0#0#�?                �C=�C=@                H�4H�4@                0#0#@        ��/����?        *���>�]@G��t��V@����]@���W@1����/C@��+��+4@���W@1����/C@��+��+@���b:P@D�JԮD1@0#0# @&�}��O@D�JԮD1@        ��#��@@��|��,@        �,����7@0����/@        ��#��0@0����/@        ���>��,@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                z�5��(@                ��#�� @�cp>@        ��#���?��/����?                ��/����?        ��#���?                ��#���?��/����?        ��#���?                        ��/����?        ���>��@                �k(��"@0����/#@        ��#�� @��/���@                ��/���@        ��#�� @                ���>��@��/����?                ��/����?        ���>��@                Lp�}>@�cp>@        ��#�� @�cp>@                �cp>@        ��#�� @                +�����;@                �k(��"@                �k(��2@                ��#���?        0#0# @                0#0# @��#���?                *�����;@鰑5@H�4H�4@��#��@���-��*@        ��#��@�cp>@        ��#�� @                ��#�� @�cp>@        ��#�� @��/����?                ��/����?        ��#�� @                        ��/����?                鰑%@                ��/����?                0����/#@        �,����7@��/���@H�4H�4@�,����7@�cp>@H�4H�4@�k(���5@�cp>@                ��/����?        �k(���5@��/����?        �k(���5@��/����?        ��#��0@                ;��,��@��/����?        ;��,��@                        ��/����?                ��/����?        ��#�� @        H�4H�4@��#�� @                                H�4H�4@        0����/@                ��/����?                �cp>@                        �A�A.@��b:��:@e#6�aJ@^��Y��X@�k(��"@On��O0@H�4H�4@z�5��@        0#0# @z�5��@                                0#0# @z�5��@On��O0@0#0#�?z�5��@0����/@0#0#�?        0����/@        z�5��@        0#0#�?��#���?        0#0#�?��#���?                                0#0#�?;��,��@                        �cp>'@                ��/����?                鰑%@        ��,���1@<l��F:B@A�s?��W@��#��0@���-��:@H�4H�4H@���>��,@��On�8@�A�A>@\Lg1��&@�cp>7@H�4H�4(@��#�� @���-��@��+��+$@��#�� @���-��@H�4H�4@        �cp>@        ��#�� @��/���@H�4H�4@��#���?                ��#���?��/���@H�4H�4@��#���?��/���@0#0#�?                0#0#�?��#���?��/���@                �cp>@        ��#���?��/����?        ��#���?                        ��/����?                        0#0# @                �C=�C=@�k(��"@On��O0@0#0# @��#�� @��/���@0#0# @��#���?��/���@0#0# @��#���?        0#0# @��#���?                                0#0# @        ��/���@        ���>��@                ��#���?��On�(@                ��/���@        ��#���?0����/@        ��#���?                        0����/@        z�5��@��/����?vb'vb'2@        ��/����?vb'vb'2@        ��/����?0#0#@        ��/����?                        0#0#@                �C=�C=,@z�5��@��/����?        ��#�� @                ��#���?��/����?                ��/����?        ��#���?                ��#�� @��/����?vb'vb'2@��#�� @��/����?vb'vb'"@��#�� @        0#0# @��#�� @                                0#0# @        ��/����?0#0#�?        ��/����?                        0#0#�?                vb'vb'"@��#���?/����/#@8k�6k�G@��#���?/����/#@��)��)3@                vb'vb'"@��#���?0����/#@��+��+$@        ��/���@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@        ��#���?��/����?vb'vb'"@��#���?��/����?0#0# @��#���?��/����?                ��/����?        ��#���?��/����?                ��/����?        ��#���?                                0#0# @                �C=�C=@                �C=�C=<@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��UhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKɅ�h��B�+         �                 ���b?���(>�?+      �����}@       �                 0��?�ޢ�e��?�       ��f$��v@       �                 P�}A?"��U�+�?�       ;��.Xt@       a                 ~`���?n��X�?�       �W��o@                          ҏ�?2��"�?j       C#mx�d@                           �?�O
�*Q�?       �͉V�M2@       
                 @��.?l�r{��?       e�6� @       	                 `F|[?f%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �               0����/@������������������������       �               鰑%@       @                 p9�? j�צ��?]       �雽�]b@       ;                 0��?
�����?>       �AC��W@                         �P��?jMg���?;       O����V@                         >�\?(���?       lz3��9@                        `r�f?f%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?                        ����?p�m ��?       �*�Ѿ6@������������������������       �               0#0#�?������������������������       �      ��       �k(���5@                          \��?�ё��?+       �w8�_P@                        �Qɰ?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?       2                 xF|�?��Yp��?'       �闭�N@       +                    �?q����?       הn�vC@       (                  L��?ڢ����?       R�T3;=;@       #                 �T?������?       Wd�R�d6@                          �~��?j��H��?       v�I�@������������������������       �               ��/����?!       "                 p���?ܗZ�	7�?       j~���@������������������������       �      �<       ��/����?������������������������       �               z�5��@$       '                 ����?k� ѽ?       �����.@%       &                 P�Zf?p����?       P	K��@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?������������������������       �      ��       ��#�� @)       *                 0i,�?���mf�?       寠�?b@������������������������       �      ��       ��/���@������������������������       �               0#0#�?,       /                 p���?��I@�?       �2d�%@-       .                  P�J�?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?0       1                 ���x?`�r{��?       e�6� @������������������������       �      ��       ���-��@������������������������       �               ��#���?3       4                    �?�v^�n�?       ��m�7@������������������������       �               ���>��,@5       :                 `x5�?fn����?       ��Y-"@6       7                  Ц6�?���/��?       @z$S��@������������������������       �               ��/����?8       9                 �^�?����?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?������������������������       �               z�5��@<       =                 P�s�?�@G���?       hu��@������������������������       �               ��/����?>       ?                  Ц6�?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?A       B                 �q�?`-�@�?       �"����I@������������������������       �               ���>��@C       \                 pִ�?�z�M�@�?       �vNF@D       Y                 `��?�?w���?       ��<��JC@E       T                 ���?�0���6�?       ���b�L@@F       I                 �$��?�u.��?       o%��z8@G       H                 �Q�?X�ih�<�?       ��
@������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?J       Q                 p���?�J	lu�?
       �a�-x1@K       P                 �n��?x���A�?       0gX\-@L       M                 p��?e��}�?       ��Se+@������������������������       �               0����/#@N       O                 �K��?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �      �<       ��#���?R       S                 �^��?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?U       X                    �?f,���O�?       ���/> @V       W                 �8�?T����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �               ��+��+@Z       [                 �/��?���/��?       @z$S��@������������������������       �               �cp>@������������������������       �               z�5��@]       `                  %��?��]ۀ��?       F���O@^       _                 ����?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?������������������������       �               ��#���?b       y                 �=jj?��q����?6       [�D�x�U@c       v                  ��d�?�2ڱ�/�?,       �ѥ|�jR@d       e                 ���#?8RL�M^�?       �)>�C@������������������������       �               �P^Cy/@f       u                 @F��hls�)�?       n+͆��7@g       p                    �?&X���`�?       �� ��4@h       i                 `�]?4=�%�?	       t=�x�-@������������������������       �               ��#��@j       m                  �G?�?R�ђ���?       �oFݜh%@k       l                  `��?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @n       o                 X/U?      �<       ��/���@������������������������       �               �cp>@������������������������       �               0����/@q       r                  �d�?ģ���c�?       �>�!J!@������������������������       �               ��/����?s       t                 l���?�zœ���?       IG���t@������������������������       �               z�5��@������������������������       �               0#0#�?������������������������       �               z�5��@w       x                 (=��>      �<       Fy�5A@������������������������       �               ��#�� @������������������������       �               ���b:@@z       {                    �?��X�?
       ���q,@������������������������       �               ��/����?|       �                 �a��?	)����?       *�GH(@}       �                  �Q�?�^h����?       S,��q$@~                        �]%�?غW�w��?       �'DQm"@������������������������       �      �<       ���>��@�       �                  E(�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               0#0#�?������������������������       �      ȼ       ��/����?�       �                 @-{V?��c�R�?2       "��S#R@�       �                  p��?$m�����?$       _d����J@�       �                 �w}�?��
��<�?"       *d�HI@�       �                 ��@�?��}g7��?       O@~a�>@�       �                 h��?      �<       /����/3@������������������������       �               �cp>@������������������������       �               On��O0@�       �                 �@�h?��F���?       :�.�-'@������������������������       �               ��#���?������������������������       �      ��       鰑%@�       �                 �3e�?4=�%�?       �(J��3@�       �                 ��y�?<9�)\e�?       _���b @�       �                ��W�y?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               ��#��@�       �                 �:��?̔fm���?       �0��z'@�       �                 ��?P�ђ���?       �oFݜh%@������������������������       �               ��#�� @�       �                 @�m�?      �<       D�JԮD!@������������������������       �               ��/����?������������������������       �               ��/���@������������������������       �      �<       ��#���?�       �                 b���?      �<       H�4H�4@������������������������       �               0#0# @������������������������       �               0#0#�?�       �                  �Q�?������?       ԋ]!_�2@������������������������       �               ��/���@�       �                  Pmj�?�Yj��}�?       ����=.@������������������������       �               ��/����?�       �                 ���?�S��W��?	       "$�
�g*@�       �                  ���?�FO���?       �ߌ$@�       �                 ؽkz?����?       ��X�)B@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?������������������������       �      ��       z�5��@�       �                 �_\�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 ��ɚ?���&�?       �S���;E@�       �                 @�l�?�J���?       ��*]Y @������������������������       �               0#0#@������������������������       �               ��#��@������������������������       �               S2%S2%A@�       �                 �6Sz?�r��-�?C       ����YZ@�       �                  �g<�?���};��?       ��;̑�5@������������������������       �               �cp>@�       �                 �L��?&�
Fq�?       /��3@�       �                 �lw?�6��b�?       &�|�1@������������������������       �      �<
       �A�A.@�       �                 �q�?x�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �      ȼ       ��/����?�       �                 @["�?p��� r�?3       ��Ģ��T@�       �                 �Sպ?��AA#�?       �>�:@������������������������       �        
       vb'vb'2@�       �                 @�ш?�~�&��?       ?�]��@������������������������       �               0#0#@�       �                 @L��?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?�       �                 �_�?{�JѠ?$       P���L@�       �                  �Ԧ�?����|e�?       �z �B�@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?�       �                 0�!�?      �<!       ������J@������������������������       �               0#0#�?������������������������       �                ��8��8J@�t�bh�hhK ��h��R�(KK�KK��h �B�  ���>��e@C�JԮDa@���Ld@���>��e@��`@B�A�P@u�}e@��`@�C=�C=<@1�����b@������S@H�4H�48@��k(/T@�]�ڕ�O@��-��-5@��#���?D�JԮD1@        ��#���?���-��@        ��#���?��/����?                ��/����?        ��#���?                        0����/@                鰑%@        �b:���S@	�cp>G@��-��-5@���b:P@���-��:@0#0#@���b:P@�e�_��7@H�4H�4@\Lg1��6@��/����?0#0#�?��#���?��/����?                ��/����?        ��#���?                �k(���5@        0#0#�?                0#0#�?�k(���5@                <��,��D@h
��6@0#0# @        �cp>@0#0#�?        �cp>@                        0#0#�?<��,��D@0����/3@0#0#�?;��,��4@On��O0@0#0#�?��,���1@D�JԮD!@0#0#�?��,���1@0����/@        z�5��@��/���@                ��/����?        z�5��@��/����?                ��/����?        z�5��@                ���>��,@��/����?        z�5��@��/����?        z�5��@                        ��/����?        ��#�� @                        ��/���@0#0#�?        ��/���@                        0#0#�?z�5��@��/���@        ��#�� @��/����?        ��#�� @                        ��/����?        ��#���?���-��@                ���-��@        ��#���?                <��,��4@�cp>@        ���>��,@                z�5��@�cp>@        z�5��@�cp>@                ��/����?        z�5��@��/����?        z�5��@                        ��/����?        z�5��@                        �cp>@0#0#�?        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?�P^Cy/@0����/3@S2%S2%1@���>��@                ��#�� @0����/3@S2%S2%1@���>��@:l��F:2@��8��8*@��#��@��/���.@��8��8*@��#�� @��/���.@�C=�C=@        ��/����?H�4H�4@                H�4H�4@        ��/����?        ��#�� @��|��,@0#0#�?��#�� @��On�(@        ��#���?��On�(@                0����/#@        ��#���?�cp>@        ��#���?                        �cp>@        ��#���?                        ��/����?0#0#�?                0#0#�?        ��/����?        ��#�� @        H�4H�4@��#�� @        0#0#�?                0#0#�?��#�� @                                ��+��+@z�5��@�cp>@                �cp>@        z�5��@                ��#���?��/����?0#0#@        ��/����?0#0#@                0#0#@        ��/����?        ��#���?                j1��tVQ@��/���.@H�4H�4@�P^CyO@鰑%@0#0#�?*�����;@鰑%@0#0#�?�P^Cy/@                z�5��(@鰑%@0#0#�?�k(��"@鰑%@0#0#�?z�5��@D�JԮD!@        ��#��@                ��#�� @D�JԮD!@        ��#�� @��/����?                ��/����?        ��#�� @                        ��/���@                �cp>@                0����/@        z�5��@��/����?0#0#�?        ��/����?        z�5��@        0#0#�?z�5��@                                0#0#�?z�5��@                Fy�5A@                ��#�� @                ���b:@@                ���>��@0����/@0#0# @        ��/����?        ���>��@�cp>@0#0# @���>��@��/����?0#0# @���>��@��/����?0#0#�?���>��@                        ��/����?0#0#�?        ��/����?                        0#0#�?                0#0#�?        ��/����?        �k(��2@��On�H@0#0#@�k(��"@�)�B�D@H�4H�4@�k(��"@�)�B�D@        ��#���?�_��e�=@                /����/3@                �cp>@                On��O0@        ��#���?鰑%@        ��#���?                        鰑%@        ��#�� @�cp>'@        ;��,��@�cp>@        ��#���?�cp>@                �cp>@        ��#���?                ��#��@                z�5��@D�JԮD!@        ��#�� @D�JԮD!@        ��#�� @                        D�JԮD!@                ��/����?                ��/���@        ��#���?                                H�4H�4@                0#0# @                0#0#�?�k(��"@D�JԮD!@0#0#�?        ��/���@        �k(��"@0����/@0#0#�?        ��/����?        �k(��"@�cp>@0#0#�?�k(��"@��/����?        z�5��@��/����?        z�5��@                        ��/����?        z�5��@                        ��/����?0#0#�?                0#0#�?        ��/����?        ��#��@        ��)��)C@��#��@        0#0#@                0#0#@��#��@                                S2%S2%A@        0����/#@C�s?��W@        �cp>@0#0#0@        �cp>@                �cp>@0#0#0@        ��/����?0#0#0@                �A�A.@        ��/����?0#0#�?                0#0#�?        ��/����?                ��/����?                ��/���@�6k�6�S@        �cp>@%S2%S27@                vb'vb'2@        �cp>@��+��+@                0#0#@        �cp>@0#0#�?        �cp>@                        0#0#�?        ��/����?�C=�C=L@        ��/����?H�4H�4@                H�4H�4@        ��/����?                        ������J@                0#0#�?                ��8��8J@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��DphFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKۅ�h��B�/         �                 ���?v�ƴ~C�?*      Ƨ�@v}@       �                  �E�?��F�z�?�       �][��w@       �                  ���?D�?��?�       _�c��r@       g                 ���?���q�?�       ��Dq@       @                 0?�pf�_�?y       �O~z�ei@       !                  �P��? ��?F       �O�էz]@                        �w�m?�Qn���?$       P��Ҵ�P@                        P�1?rF9i5�?       j�HhH9@	       
                  �"�?��|��?       ���ĺw@������������������������       �      ��       ��/���@                        lS�a?Zn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @                         <�e?`n����?       ��Y-2@                        @Ws�?�d�$���?       <��#�.@                        �r��?@9�)\e�?       _���b @������������������������       �               ;��,��@������������������������       �               �cp>@������������������������       �      ��       ���>��@                        �ori?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?                        ��ͅ?4K����?       j�TqŏD@                         T�u?x7uV��?       m}�'�:@                         p��?��6L�n�?       �E#��h @������������������������       �               ��/����?������������������������       �      �<       ���>��@������������������������       �        
       �k(��2@                         ��Ӈ?$�b���?       �GXvƒ,@                        ��ʵ?|�G���?       ��%�|@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               ;��,��$@"       7                 �'�l?�tȠ�,�?"       �xC��I@#       0                  �6�?�[ޞ�?       �N�m?@$       /                 �mEr?�y�8��?
       87@�-@%       .                 ���뾺�k{��?	       `;�W� *@&       -                 P#%v?f%@�"�?       �6�E�!@'       (                   \��?Ɣfm���?       ��Z�N@������������������������       �               0����/@)       *                 �}#$?\n����?       � ��w<@������������������������       �               ��#���?+       ,                 `�)Q?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#���?������������������������       �               ��#��@������������������������       �      м       ��/����?1       2                 �#�t?bsfi��?	       3��w�0@������������������������       �               ��/���@3       4                 �4?�����?       �v�qp�!@������������������������       �               H�4H�4@5       6                 x��?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �               0����/@8       ;                 �j��?����?       8�nN�R4@9       :                 ��͑?Xb8�Y�?	       HJͰ(@������������������������       �      �<       \Lg1��&@������������������������       �      ȼ       ��/����?<       =                 ����?���/��?       U��7�@������������������������       �               z�5��@>       ?                  Ц6�?$ k�Lj�?       �q��l}@������������������������       �      �<       ��/���@������������������������       �               ��#���?A       b                 p�3g?����?3       ;O?QU@B       ]                  ��d�?Dg3E��?,       �o��FWR@C       F                  �X?]\��?(       G��(JP@D       E                 @�Ks?���/��?       @z$S��@������������������������       �               �cp>@������������������������       �               z�5��@G       L                  �`�?/�W�>�?%       E�it�M@H       I                 @F��pP'�'�?       B�nm��?@������������������������       �               �cp>7@J       K                    �?)���?       y��uk!@������������������������       �               ��/���@������������������������       �               ��#���?M       T                  @mj�?J%?�)�?       C?�e�p;@N       O                  ��?��%�U��?       o/o�a2@������������������������       �               ��#���?P       S                 �6�?������?       �N0gX1@Q       R                 @�i�?�`@s'��?       Ei_y,*@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �      �<       鰑%@U       \                 �^1�?H��aB��?       ����"@V       W                 �F��?����]L�?       N66�ͯ@������������������������       �               ��#���?X       Y                  �P�?�@G���?       hu��@������������������������       �               0#0#�?Z       [                 pU�<?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��#��@^       _                 ���?��6L�n�?       �E#��h @������������������������       �               ;��,��@`       a                 ��T?bn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @c       d                 �+�[?h��`p��?       �����'@������������������������       �               �cp>@e       f                   ��?X*�'=P�?        �2"@������������������������       �               ��/����?������������������������       �               0#0# @h       y                 `���?.F%?��?-       RS)AQ@i       r                 ��)�?w`��?       � �D@j       o                 �;�?j�а.�?       ��W�&2@k       l                 �ʌ�?���Ww�?	       x��4]�,@������������������������       �               ZLg1��&@m       n                8�/��?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?p       q                pT�?      �<       ��/���@������������������������       �               �cp>@������������������������       �               ��/����?s       t                 �$I�?(��*ʽ�?       	�t�U7@������������������������       �               �cp>@u       x                 P�u�?��[\��?       )sh�24@v       w                 ���?�o���?       o�9�F@������������������������       �               0#0#@������������������������       �               ��#���?������������������������       �        	       �A�A.@z       {                 P�Ƥ?f��o�3�?       J<��;@������������������������       �               �k(��"@|       }                 ��?�qL�Ľ�?       <W�w�y2@������������������������       �               ��/����?~                        ��?��G�MJ�?       F�v�Q�1@������������������������       �               z�5��@�       �                 @�	�?���BK�?	       �)��؜&@�       �                 `m�?�J���?       a���@�       �                 ��s'?�zœ���?       IG���t@������������������������       �               0#0#�?������������������������       �               z�5��@������������������������       �               0#0# @������������������������       �      �<       ;��,��@�       �                 `���?�ld���?       ���$]Z:@�       �                  v��?���_`�?       &!j�\+"@�       �                 �'��?�26�
�?       4��*8E@�       �                 �z?�djH�E�?       ^�\m�n@������������������������       �               ��#��@�       �                 �h�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ȼ       ��/����?������������������������       �               0#0# @������������������������       �               E�JԮD1@�       �                 �6SZ?YtT_��?<       Sb�ۙ�T@�       �                 �Y`�?��B�rM�?'       �"�͑vK@�       �                 ���@?Ȫ�a��?#       ��h6iH@�       �                 h'x�?VƲ�<|�?       !�[�C@�       �                 ��n?�f%j��?       ��ꁞ9<@�       �                  ��>l@ȱ��?       nm���S@������������������������       �               ��#���?������������������������       �      ��       0����/@�       �                  5��?������?       Xd�R�d6@�       �                 �-�?#����?       x�߄�3@������������������������       �               ��/����?�       �                  p�:?�hK)�?       �h��K�2@������������������������       �      ��	       ���>��,@�       �                 p#��?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@�       �                 (��u?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?�       �                 �/��?��_~"��?       �bj��%@������������������������       �               �cp>@�       �                 ��½?@��X�&�?       �6��	�@������������������������       �               ��/����?�       �                 𝠬?£���c�?       �>�!J!@������������������������       �               z�5��@�       �                    �?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                  2�M?���k�L�?       sk��#@������������������������       �               �cp>@�       �                  ��M�?�3`���?       .�r��@�       �                 �f�V?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               0#0# @�       �                 ����?�D#���?       �B�j@������������������������       �               0#0#@������������������������       �               ��#�� @�       �                 0�]Z?      �<       �C=�C=<@������������������������       �               0#0#�?������������������������       �               �;�;;@�       �                 p��z?�sU���?:       V�*e�jV@�       �                 @Mί?��O����?'       Ԧ���7O@�       �                  ��?��yO�?       �a)5':@�       �                 �Ҕ?e��}�?       ��Se+@������������������������       �               ��#���?������������������������       �               ��On�(@�       �                  \��?Ħ54�3�?       W���)@�       �                 �{�?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 0vb�?�?�0�!�?       a`�T�$@������������������������       �               vb'vb'"@������������������������       �      ȼ       ��/����?�       �                   ��?T�/J�?       ��"Wg�A@�       �                  �Mm�?���9��?       l�P"��)@�       �                  �!�?�@G���?       hu��@�       �                 ���?|�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               ��/���@������������������������       �               ��+��+@�       �                 `�1�? ��:y�?       7��7@�       �                 �c�?ȏ�yŷ?       L�j>�45@�       �                 ���?�D#���?       �B�j@������������������������       �               0#0#�?�       �                  X��?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               vb'vb'2@������������������������       �      ȼ       ��/����?�       �                  p�{�?      �<       �;�;;@������������������������       �               0#0#�?������������������������       �               ��8��8:@�t�bh�hhK ��h��R�(KK�KK��h �B�  �>��d@�H��tXe@bF`�a@������c@��z��wb@��)��)S@��#��`@*����-_@�ڬ�ڬD@���b:`@`#6�aZ@��)��)C@���W@�e�_��W@�A�A.@��Gp_R@2����/C@H�4H�4@�}�\I@���-��*@0#0# @���>��,@鰑%@        ��#�� @0����/@                ��/���@        ��#�� @��/����?                ��/����?        ��#�� @                z�5��(@�cp>@        z�5��(@�cp>@        ;��,��@�cp>@        ;��,��@                        �cp>@        ���>��@                        �cp>@                ��/����?                ��/����?        �YLg1B@�cp>@0#0# @�#���9@��/����?        ���>��@��/����?                ��/����?        ���>��@                �k(��2@                <��,��$@��/����?0#0# @        ��/����?0#0# @                0#0# @        ��/����?        ;��,��$@                \Lg1��6@��On�8@0#0#@���>��@&jW�v%4@0#0#@���>��@��/���@        ���>��@�cp>@        z�5��@�cp>@        ��#�� @�cp>@                0����/@        ��#�� @��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                ��#���?                ��#��@                        ��/����?                ��On�(@0#0#@        ��/���@                0����/@0#0#@                H�4H�4@        0����/@0#0#�?                0#0#�?        0����/@        �P^Cy/@0����/@        \Lg1��&@��/����?        \Lg1��&@                        ��/����?        ��#��@��/���@        z�5��@                ��#���?��/���@                ��/���@        ��#���?                �k(��2@��|��L@vb'vb'"@�k(��2@���-��J@0#0#�?ZLg1��&@c#6�aJ@0#0#�?z�5��@�cp>@                �cp>@        z�5��@                ��#�� @��On�H@0#0#�?��#���?��/���>@                �cp>7@        ��#���?��/���@                ��/���@        ��#���?                ���>��@0����/3@0#0#�?��#�� @Nn��O0@        ��#���?                ��#���?On��O0@        ��#���?�cp>@                �cp>@        ��#���?                        鰑%@        ;��,��@�cp>@0#0#�?��#���?�cp>@0#0#�?��#���?                        �cp>@0#0#�?                0#0#�?        �cp>@                ��/����?                ��/����?        ��#��@                ���>��@��/����?        ;��,��@                ��#�� @��/����?                ��/����?        ��#�� @                        ��/���@0#0# @        �cp>@                ��/����?0#0# @        ��/����?                        0#0# @�YLg1B@0����/#@%S2%S27@z�5��(@D�JԮD!@��+��+4@[Lg1��&@�cp>@0#0#�?\Lg1��&@��/����?0#0#�?ZLg1��&@                        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/���@                �cp>@                ��/����?        ��#���?�cp>@��)��)3@        �cp>@        ��#���?        ��)��)3@��#���?        0#0#@                0#0#@��#���?                                �A�A.@�,����7@��/����?H�4H�4@�k(��"@                ���>��,@��/����?H�4H�4@        ��/����?        ���>��,@        H�4H�4@z�5��@                ��#�� @        H�4H�4@z�5��@        H�4H�4@z�5��@        0#0#�?                0#0#�?z�5��@                                0#0# @;��,��@                ��#��@1����/3@H�4H�4@��#��@��/����?H�4H�4@��#��@��/����?0#0#�?��#��@��/����?0#0#�?��#��@                        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?                        0#0# @        E�JԮD1@        |�5��8@�cp>7@eJ�dJ�A@|�5��8@�cp>7@�C=�C=@\Lg1��6@�cp>7@H�4H�4@�k(���5@Nn��O0@0#0#�?�k(��2@/����/#@        ��#���?0����/@        ��#���?                        0����/@        ��,���1@0����/@        ��,���1@��/����?                ��/����?        ��,���1@��/����?        ���>��,@                z�5��@��/����?                ��/����?        z�5��@                        �cp>@                ��/����?                ��/����?        z�5��@���-��@0#0#�?        �cp>@        z�5��@��/���@0#0#�?        ��/����?        z�5��@��/����?0#0#�?z�5��@                        ��/����?0#0#�?                0#0#�?        ��/����?        ��#���?���-��@0#0# @        �cp>@        ��#���?��/����?0#0# @��#���?��/����?        ��#���?                        ��/����?                        0#0# @��#�� @        0#0#@                0#0#@��#�� @                                �C=�C=<@                0#0#�?                �;�;;@z�5��@�cp>7@Q��N��O@z�5��@�cp>7@xb'vb'B@��#�� @��/���.@vb'vb'"@��#���?��On�(@        ��#���?                        ��On�(@        ��#���?�cp>@vb'vb'"@��#���?��/����?        ��#���?                        ��/����?                ��/����?vb'vb'"@                vb'vb'"@        ��/����?        ��#���?��/���@�;�;;@        �cp>@�C=�C=@        �cp>@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @        ��/���@                        ��+��+@��#���?��/����?��+��+4@��#���?        ��+��+4@��#���?        0#0# @                0#0#�?��#���?        0#0#�?                0#0#�?��#���?                                vb'vb'2@        ��/����?                        �;�;;@                0#0#�?                ��8��8:@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ%�[6hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKۅ�h��B�/         �                 ��ז?֙�M�?-      ��̚щ}@       w                 ��?_�D���?�       3�i�̅u@                        ���W?�=[|�{�?�       s/�tm@                        � �l?�&��$C�?       ���+p8@       
                 ���2?���.�2�?       ��k	j3@                        ��g�?l��H��?       v�I�@������������������������       �               ��#�� @       	                 ��E?& k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?������������������������       �      �<
       ��On�(@                         \��?�Z�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@                          ҏ�?h�x���?�       ~i��fj@                        |ίd?��Xv#�?       (RҀh�4@                        ૗l?��Z�	7�?       j~���@������������������������       �               z�5��@������������������������       �      �<       ��/����?                        �?p�r{��?       e�6� /@������������������������       �               ��#���?                          �g�?��&���?       ��G2��,@������������������������       �               ��/���@                        ��k�?�`@s'��?       Fi_y,*@                        �U�,?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?                           �?      �<       ��/���@������������������������       �               ��/����?������������������������       �               ��/����?       (                  1�>"Rz�O��?u       :���g@        !                 ��{?.�~�!�?       Lƿ�;q*@������������������������       �               ;��,��@"       '                  @���?r^�(���?       � K�h @#       &                 @��?`�ih�<�?       ��
@$       %                 (�i<?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               0#0#@������������������������       �               ��#���?)       Z                 ���O?�b<ʚ��?n       �"ͯ.f@*       =                 �Ӻs?dZ����?I       R�VȎ^@+       <                 �G�? �`�k	�?)       �-�y�Q@,       /                  �Q�?�����?       9�nN�RD@-       .                 3Ё$?f%@�"�?       ��[�@������������������������       �      �<       ��/���@������������������������       �               ��#�� @0       7                 ����?�q���?       ��|�^A@1       6                 �Y��?�]���?       �j0�W�<@2       3                 p�;?4Bms�?       ��֖��;@������������������������       �      ȼ       
�#���9@4       5                  �Q�?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �      �<       ��/����?8       ;                 �4�r?���/��?       @z$S��@9       :                  P�"�?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?������������������������       �               Jp�}>@>       W                 ��\�?���b�j�?        FgW~��I@?       @                 `s5�?���؜��?       �[u��E@������������������������       �               0#0# @A       V                 ���?��h�Z�?       �YR�D@B       C                  �\�?������?       ��W/O�C@������������������������       �               ;��,��@D       S                 �E�?�P��=.�?       ZS�i�	A@E       L                    �?�PЈ��?       U�{�>@F       G                 �h�?@H�,.̷?       �J�$r.5@������������������������       �               �cp>'@H       K                  L��?ܜ�x�?       d��إV#@I       J                 �5�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       ��/���@M       N                  �f?���1n�?       <���4�!@������������������������       �               ��#�� @O       P                 �J��?��n��?       �-H�\@������������������������       �               ��#���?Q       R                 ����?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �               0����/@T       U                 �2OF?����|e�?       �z �B�@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?������������������������       �               0#0# @X       Y                 ���?      �<       ��#�� @������������������������       �               ��#��@������������������������       �               ��#��@[       \                 ���`? f�r��?%       ����.�K@������������������������       �               ��/����?]       v                 0)��?����-��?$       0	R�b"K@^       k                 �U�?�ڹ����?#       ��}J�J@_       h                 �;�?�|]��e�?       ��Ҩ�B@`       a                 ��R?b�d����?	       4K}@0�*@������������������������       �               0#0# @b       g                 �ͪ�?2��/��?       ��t�o�&@c       f                 `��b?D�k����?       b*pn�$@d       e                 ����?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �               0#0#�?i       j                    �?      �<       [Lg1��6@������������������������       �        
       �P^Cy/@������������������������       �               ���>��@l       m                  s��?Y�Z%x
�?       C���_#1@������������������������       �               ��/���@n       q                 ����?&g���?
       ��+���*@o       p                 D2²?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @r       s                  ���?8�k����?       b*pn�$@������������������������       �               ���>��@t       u                  y��?R����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?������������������������       �     ��<       0#0#�?x       �                 �QT�?��8D�_�?B       �H�.[@y       �                 ��?hzmi0o�?:       tQ?GF%W@z                        аs}?��v�@��?0       �6��S@{       ~                 @�Dv?���o�:�?       ����+@|       }                 `A�t?r@ȱ��?       om���S@������������������������       �               0����/@������������������������       �               ��#���?������������������������       �               0#0# @�       �                 �a�?ƽ'	�_�?*       �3�R�EO@������������������������       �               0����/#@�       �                 �I�?��X�"��?"       θ%��yJ@�       �                 `�;�?�2|�?        >��#�pI@�       �                 -��?�%E�N��?       �h���2@������������������������       �               0#0#@�       �                 ���?Ђ�O���?
       �O�
|-@�       �                  `%+�?�O-r��?       �.w��e)@�       �                 �޲�?      �<       ���-��@������������������������       �               ��/����?������������������������       �               �cp>@�       �                  Fn�?���/��?       @z$S��@������������������������       �               �cp>@������������������������       �               z�5��@�       �                 ��N�? �J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?�       �                 0��?-�����?       �#$w@@�       �                 ���?�1A�]�?       ]g	��?@�       �                  �?�AP�9��?       i��6��@������������������������       �               ��+��+@������������������������       �      �<       ��/����?�       �                 x�'�?tD R�?       �xK&�8@�       �                 ��o�?      �<       E�JԮD1@������������������������       �               ��/����?������������������������       �               On��O0@�       �                  ��?��n��?       �-H�\@�       �                 �η�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               0����/@������������������������       �      �<       ��#���?�       �                  ���?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?�       �                   �P�?      �<
       0#0#0@������������������������       �               0#0# @������������������������       �        	       �C=�C=,@�       �                 �a�?      �<       0#0#0@������������������������       �               0#0# @������������������������       �               �C=�C=,@�       �                 ��?��/���?T       eƺ	`@�       �                 �Y�?|��j�?       p$��Y5@�       �                   B�?x�w�o�?
       �c/�P1@�       �                  ��^�?(Й����?	       �3�N0@�       �                 -��?��oR��?       l�Q6�(@�       �                 2>��?��q�R�?       C}Ԥ@������������������������       �               ��#���?�       �                 ��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       �k(��"@�       �                 ���?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �               0#0#@�       �                  �?�俿3�?G       ��Ʀ�Z@�       �                 @=��?���mf�?       寠�?b@������������������������       �      ��       ��/���@������������������������       �               0#0#�?�       �                 0��?8��G��?C       ��΂�Y@�       �                 pJ�q?�V����?7       �i�96:U@�       �                  `ۣ?��?�5�?       0����E@�       �                 0ys8?(��`�?
       П@��.(@������������������������       �               ��#��@�       �                  ��?C��X�&�?       �6��	�@�       �                 ȶI�?�zœ���?       IG���t@������������������������       �               0#0#�?������������������������       �               z�5��@������������������������       �      ��       ��/���@�       �                 Z&�?N���?       v�ܲw?@������������������������       �               �cp>@�       �                    �?���)�?       ��@#�9@�       �                 `���?l@ȱ��?       nm���S@�       �                 `TF�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ��       ��/���@�       �                 ����?����	�?       WK0�3@������������������������       �               �cp>@�       �                  Pmj�?�~�nE�?	       v��Bh 1@�       �                 @?�� ��?       rp� k@������������������������       �               0#0# @������������������������       �      �<       ��/���@�       �                  X��?r��R[�?       ��"PK&@������������������������       �               0#0# @�       �                  �6�?T����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �               �ڬ�ڬD@������������������������       �               S2%S2%1@�t�bh�hhK ��h��R�(KK�KK��h �B�  ���#8e@q�'�x�b@�i��b@��Gp_b@h>�c�^@���~�gR@YUUUU5a@r�'�x�R@#0#06@z�5��@9l��F:2@        z�5��@On��O0@        z�5��@��/���@        ��#�� @                ��#���?��/���@                ��/���@        ��#���?                        ��On�(@        z�5��@��/����?                ��/����?        z�5��@                �,���n`@��|��L@#0#06@;��,��@��/���.@        z�5��@��/����?        z�5��@                        ��/����?        ��#�� @���-��*@        ��#���?                ��#���?���-��*@                ��/���@        ��#���?�cp>@        ��#���?��/����?        ��#���?                        ��/����?                ��/���@                ��/����?                ��/����?        &�}��_@鰑E@#0#06@z�5��@��/����?H�4H�4@;��,��@                ��#���?��/����?H�4H�4@        ��/����?H�4H�4@        ��/����?0#0# @        ��/����?                        0#0# @                0#0#@��#���?                Mp�}^@�)�B�D@0#0#0@������S@����z�A@0#0# @��>���N@/����/#@        �P^Cy?@0����/#@        ��#�� @��/���@                ��/���@        ��#�� @                ���>��<@�cp>@        �#���9@�cp>@        �#���9@��/����?        
�#���9@                        ��/����?                ��/����?                ��/����?                ��/����?        z�5��@�cp>@        z�5��@��/����?                ��/����?        z�5��@                        ��/����?        Jp�}>@                ��,���1@�cp>�9@0#0# @�k(��"@�cp>�9@0#0# @                0#0# @�k(��"@�cp>�9@H�4H�4@�k(��"@�cp>�9@0#0#@;��,��@                ��#��@�cp>�9@0#0#@��#��@��On�8@0#0#�?��#���?'jW�v%4@                �cp>'@        ��#���?E�JԮD!@        ��#���?��/����?                ��/����?        ��#���?                        ��/���@        z�5��@0����/@0#0#�?��#�� @                ��#���?0����/@0#0#�?��#���?                        0����/@0#0#�?                0#0#�?        0����/@                ��/����?H�4H�4@                H�4H�4@        ��/����?                        0#0# @��#�� @                ��#��@                ��#��@                =��,��D@�cp>@0#0# @        ��/����?        =��,��D@0����/@0#0# @=��,��D@0����/@�C=�C=@���b:@@        0#0#@�k(��"@        0#0#@                0#0# @�k(��"@        0#0# @�k(��"@        0#0#�?��#���?        0#0#�?��#���?                                0#0#�?��#�� @                                0#0#�?[Lg1��6@                �P^Cy/@                ���>��@                �k(��"@0����/@H�4H�4@        ��/���@        �k(��"@��/����?H�4H�4@        ��/����?0#0# @        ��/����?                        0#0# @�k(��"@        0#0#�?���>��@                ��#�� @        0#0#�?��#�� @                                0#0#�?                0#0#�?�k(��"@�e�_��G@~˷|˷I@�k(��"@�e�_��G@dJ�dJ�A@�k(��"@ f�_��G@��)��)3@��#���?0����/@0#0# @��#���?0����/@                0����/@        ��#���?                                0#0# @��#�� @��]�ڕE@#0#0&@        0����/#@        ��#�� @�-����@@#0#0&@z�5��@�-����@@#0#0&@��#��@/����/#@��+��+@                0#0#@��#��@/����/#@0#0#�?z�5��@/����/#@                ���-��@                ��/����?                �cp>@        z�5��@�cp>@                �cp>@        z�5��@                ��#���?        0#0#�?                0#0#�?��#���?                ��#�� @�e�_��7@H�4H�4@��#���?�e�_��7@H�4H�4@        ��/����?��+��+@                ��+��+@        ��/����?        ��#���?h
��6@0#0#�?        E�JԮD1@                ��/����?                On��O0@        ��#���?0����/@0#0#�?��#���?        0#0#�?��#���?                                0#0#�?        0����/@        ��#���?                ��#�� @                ��#���?                ��#���?                                0#0#0@                0#0# @                �C=�C=,@                0#0#0@                0#0# @                �C=�C=,@\Lg1��6@�a#6�;@��jS@z�5��(@�cp>@H�4H�4@z�5��(@�cp>@0#0# @z�5��(@�cp>@0#0#�?;��,��$@��/����?0#0#�?��#���?��/����?0#0#�?��#���?                        ��/����?0#0#�?        ��/����?                        0#0#�?�k(��"@                ��#�� @��/����?        ��#�� @                        ��/����?                        0#0#�?                0#0#@<��,��$@��On�8@p�fm��Q@        ��/���@0#0#�?        ��/���@                        0#0#�?<��,��$@鰑5@gJ�dJ�Q@<��,��$@鰑5@������J@<��,��$@鰑5@H�4H�4(@���>��@��/���@0#0#�?��#��@                z�5��@��/���@0#0#�?z�5��@        0#0#�?                0#0#�?z�5��@                        ��/���@        z�5��@D�JԮD1@#0#0&@        �cp>@        z�5��@�cp>'@#0#0&@��#���?0����/@        ��#���?��/����?        ��#���?                        ��/����?                ��/���@        ��#�� @���-��@#0#0&@        �cp>@        ��#�� @��/���@#0#0&@        ��/���@0#0# @                0#0# @        ��/���@        ��#�� @        vb'vb'"@                0#0# @��#�� @        0#0#�?                0#0#�?��#�� @                                �ڬ�ڬD@                S2%S2%1@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�	3 hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK녔h��Bh3         �                 �0Md?���G�?)      %��L�}@       �                 �j�?��#��?�       Ρ���v@       f                 P�)�?>���[�?�       c$W��it@       a                 кI�?�`�\��?|       hJ8Ѹh@       B                 ��??riHsy��?u       �/���>f@       )                 83<p?�ۧ�`�?W       ��y�C`@                        "?��+����?8       $��IU@       	                 ~W�>�(1k��?       �ꁞ9�6@������������������������       �               ��b:��*@
                          �?`�j���?       ���z"@������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?                        P�1?
S��/��?*       �Rm�v�N@������������������������       �               ��/����?       &                 ��]"?�ө@h�?(       �����M@                         `s�?P�];�?       ��t�HA@������������������������       �               �cp>@       #                 �m��?$1_#�?       R!�M<@                         0��j?�T`�[k�?       n��F:l9@                        @.��>�)z� ��?
       ~�\�,@������������������������       �               ��#�� @                        @F����/��?	       ?z$S��'@                         ���?:ǵ3���?       �q�ͨ�@                        �C[?ޗZ�	7�?       j~���@                        @Ws�?f%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �      ��       �cp>@                        `%�7?����?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?!       "                 �'�U?      �<       ZLg1��&@������������������������       �               ��#�� @������������������������       �               �k(��"@$       %                    �?     ��<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?'       (                  `S��?���OT�?       q�>%,�9@������������������������       �               {�5��8@������������������������       �      �<       ��/����?*       ?                 ��?� ^�D��?       8 >��F@+       8                 �
o?���/��?       8��o��C@,       5                 `��T? �Ұ��?       �1��<@-       .                 ��Y?� ^�D��?       8 >��6@������������������������       �               ���-��@/       0                  �P��?:9�)\e�?       _���b0@������������������������       �               ���>��@1       4                 �5W�?b%@�"�?       �6�E�!@2       3                 ��{�?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@������������������������       �      ��       0����/@6       7                 ���?      �<       �cp>@������������������������       �               ��/����?������������������������       �               0����/@9       <                 _%?����X��?       (��֞&@:       ;                 ��p?      �<       �k(��"@������������������������       �               ��#���?������������������������       �               ��#�� @=       >                 �j��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?@       A                 (�I�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               0����/@C       X                 p��?`?2�6�?       R?���G@D       U                 0!�?N��Y�?       >�&�D@E       J                 ���@?��fƲ��?       �u�:?@F       I                 t�@`?����?       ��X�)B@G       H                  P�"�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#�� @K       R                 P�+�?�`@s'��?       Ei_y,*;@L       Q                 p6!�?|��� �?       0)���"8@M       P                 ��vi?�B�� �?       �HI�7@N       O                 �=E? ܜ�x�?       d��إV#@������������������������       �               ��#���?������������������������       �               E�JԮD!@������������������������       �               ���-��*@������������������������       �      �<       ��#���?S       T                 >�ht?Tn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @V       W                 ���N?      �<       鰑%@������������������������       �               �cp>@������������������������       �               0����/@Y       `                 �/��?bn����?       � ��w<@Z       ]                  %�r?�d�$���?       �T�f@[       \                h8�YT?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ��#�� @^       _                 h�B?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ȼ       ��/����?b       e                   ��?x��Ww�?       v��4]�,@c       d                 <�Й?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?������������������������       �               [Lg1��&@g       n                 `|)�?����ř�?T       h�u!�`@h       m                 � ��?��^���?       ���w!@i       j                 ����?xLU���?       h�ҹ^�@������������������������       �               0����/@k       l                �E9�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0#�?o       �                 �p�?g��-V�?N       �F�N@g_@p       �                      �૽���?       ԤAc�xE@q       �                 �N��?�3J��;�?       2�W�@@r       �                 P8��?H������?       m���{"9@s       |                 ��~?v쾰3�?       .=����4@t       u                 0=�?o .A��?       �wPq�/@������������������������       �               0����/@v       w                 H��?�(^:�w�?       Z�� 2&@������������������������       �               H�4H�4@x       {                 ���?ҟ��X�?       l�n�/@y       z                 x��?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               0#0# @}       �                  �Ǥ?�d�$���?       �T�f@~                        ����?      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@������������������������       �      ȼ       ��/����?������������������������       �               ��#��@������������������������       �               �C=�C=@�       �                ���v?�}/W�?	       �r�.�%@������������������������       �               0#0# @�       �                 @���?��^���?       ���w!@�       �                 pM�D?xLU���?       i�ҹ^�@�       �                    �?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �               0����/@������������������������       �               0#0#�?�       �                 0*tC?�4���?2       (t�ӪT@�       �                 PC�?��n?�?&       !z��k9P@�       �                   ��?���N���?       �-\BmC@�       �                p�qz�?2�c3���?       �uk��!@������������������������       �               ��/���@�       �                 ��{�?�d�$���?       �T�f@������������������������       �               ��#�� @�       �                 �)��?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?�       �                 `U�?a	._�?       B^��N�=@�       �                 NK�X?�}O:�ӱ?       ��d]��;@������������������������       �               0#0#�?������������������������       �               ��b:��:@�       �                 ���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 ���?t��7��?       6��u{:@������������������������       �               �cp>@�       �                  pjS�?���)��?       T���*7@�       �                 `�x�?���N���?       �O��!3@�       �                  ��?��b�}�?       �1%
�-@�       �                  �[??�|2N��?       �3K}@������������������������       �               z�5��@������������������������       �               0#0# @�       �                 ���?ZV�IS��?       '���d�#@�       �                  ���?���/��?       @z$S��@������������������������       �      ��       z�5��@�       �                 @*��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?�       �                  `�J�?�@G���?       hu��@������������������������       �               0#0#�?�       �                 艝�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �               0#0#@�       �                  /�u?Q�aɴ�?       �Sy��1@������������������������       �               �cp>@�       �                 `w9�?Ǔ�R �?       ��u�(@������������������������       �               z�5��@�       �                    �?�֪u�_�?       ��?�8@������������������������       �               ��/���@�       �                   �x�?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 ��˺?6���t�?       mMU2 �A@������������������������       �               ��/���@�       �                 �xѱ?,!�IPD�?       �O�S�
@@�       �                 Фͽ?��Dr�?       �9[�7�!@������������������������       �               ��/����?�       �                pn�ǣ?���1p8�?       |곯�@�       �                 0I��?�@����?       ���a�@�       �                  ���?z��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               0#0# @�       �                   .p�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                  �?z�&�?       �ۄ-7@�       �                 �qg�?�*����?       �=��76@�       �                 �D;�?7��b�?	       %�|�1@�       �                 �G\�?X�ih�<�?       ��
@������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?������������������������       �      ��       ��+��+$@�       �                 p�h�?�|2N��?       �3K}@������������������������       �               z�5��@������������������������       �               0#0# @������������������������       �      �<       ��/����?�       �                 Pt%�?p>�0�!�?D       �D�4��[@�       �                 P�!z?�AP�9��?       h��6��+@������������������������       �               vb'vb'"@�       �                 ��3�?���mf�?       寠�?b@�       �                ��ϖ�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       �cp>@�       �                 ��W�?��]�@��?<       <M��xX@�       �                  �E�?�՜���?&       �
�#�N@�       �                  ���?�n���k�?       4��&�:@������������������������       �               H�4H�48@�       �                 xs�?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �      м       dJ�dJ�A@�       �                  ���?T�ih�<�?       s���͆A@������������������������       �               �cp>@�       �                 p1m�?(r����?       Qz�i@@������������������������       �      ��       k�6k�69@�       �                 v�2�?�AP�9��?       i��6��@������������������������       �               ��/����?������������������������       �               ��+��+@�t�b��&     h�hhK ��h��R�(KK�KK��h �B  ���>��e@����Xb@��)��)c@���>��e@��t�Ha@������J@u�}e@�]�ڕ�_@=�C=�C?@�>��n[@��-��bT@0#0#�?ZUUUU�X@g
���S@        �k(���U@��]�ڕE@        ��#��P@:l��F:2@        �k(���5@��/����?        ��b:��*@                ��#�� @��/����?        ��#�� @                        ��/����?        �GpAF@D�JԮD1@                ��/����?        �GpAF@��/���.@        ������3@��|��,@                �cp>@        ������3@D�JԮD!@        ������3@�cp>@        ��#�� @�cp>@        ��#�� @                z�5��@�cp>@        z�5��@0����/@        z�5��@��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#�� @                        �cp>@        z�5��@��/����?        z�5��@                        ��/����?        ZLg1��&@                ��#�� @                �k(��"@                        �cp>@                ��/����?                ��/����?        {�5��8@��/����?        {�5��8@                        ��/����?        <��,��4@��On�8@        ;��,��4@0����/3@        <��,��$@:l��F:2@        <��,��$@��On�(@                ���-��@        <��,��$@�cp>@        ���>��@                z�5��@�cp>@        z�5��@��/����?                ��/����?        z�5��@                        0����/@                �cp>@                ��/����?                0����/@        <��,��$@��/����?        �k(��"@                ��#���?                ��#�� @                ��#���?��/����?        ��#���?                        ��/����?                �cp>@                ��/����?                0����/@        ZLg1��&@:l��F:B@        ���>��@E�JԮDA@        ���>��@�e�_��7@        z�5��@��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#�� @                ��#��@�cp>7@        ��#�� @h
��6@        ��#���?h
��6@        ��#���?D�JԮD!@        ��#���?                        E�JԮD!@                ���-��*@        ��#���?                ��#�� @��/����?                ��/����?        ��#�� @                        鰑%@                �cp>@                0����/@        ��#��@��/����?        ��#��@��/����?        z�5��@                ��#���?                ��#�� @                ��#���?��/����?                ��/����?        ��#���?                        ��/����?        ZLg1��&@��/����?0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?[Lg1��&@                    �M@�'�xr�F@�A�A>@        ���-��@0#0# @        ���-��@0#0#�?        0����/@                ��/����?0#0#�?                0#0#�?        ��/����?                        0#0#�?    �M@2����/C@�C=�C=<@;��,��$@���-��*@��)��)3@;��,��$@���-��@�A�A.@;��,��$@���-��@0#0# @z�5��@���-��@0#0# @��#�� @�cp>@0#0# @        0����/@        ��#�� @��/����?0#0# @                H�4H�4@��#�� @��/����?0#0# @��#�� @��/����?                ��/����?        ��#�� @                                0#0# @��#��@��/����?        ��#��@                ��#���?                z�5��@                        ��/����?        ��#��@                                �C=�C=@        ���-��@0#0#@                0#0# @        ���-��@0#0# @        ���-��@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        0����/@                        0#0#�?4��tSH@��On�8@vb'vb'"@���#8E@��|��,@0#0# @���b:@@�cp>@0#0#�?��#��@0����/@                ��/���@        ��#��@��/����?        ��#�� @                ��#�� @��/����?        ��#�� @                        ��/����?        *�����;@��/����?0#0#�?��b:��:@        0#0#�?                0#0#�?��b:��:@                ��#���?��/����?                ��/����?        ��#���?                <��,��$@D�JԮD!@�C=�C=@        �cp>@        ;��,��$@�cp>@�C=�C=@;��,��$@�cp>@H�4H�4@z�5��@�cp>@H�4H�4@z�5��@        0#0# @z�5��@                                0#0# @z�5��@�cp>@0#0#�?z�5��@�cp>@        z�5��@                        �cp>@                ��/����?                ��/����?                �cp>@0#0#�?                0#0#�?        �cp>@                ��/����?                ��/����?        ��#��@                                0#0#@z�5��@鰑%@0#0#�?        �cp>@        z�5��@0����/@0#0#�?z�5��@                        0����/@0#0#�?        ��/���@                ��/����?0#0#�?        ��/����?                        0#0#�?��#��@/����/#@#0#06@        ��/���@        ��#��@�cp>@#0#06@��#���?��/���@0#0#@        ��/����?        ��#���?��/����?0#0#@        ��/����?0#0#@        ��/����?0#0# @                0#0# @        ��/����?                        0#0# @��#���?��/����?                ��/����?        ��#���?                z�5��@��/����?vb'vb'2@z�5��@��/����?vb'vb'2@        ��/����?0#0#0@        ��/����?H�4H�4@                H�4H�4@        ��/����?                        ��+��+$@z�5��@        0#0# @z�5��@                                0#0# @        ��/����?                鰑%@g'vb'�X@        ��/���@��+��+$@                vb'vb'"@        ��/���@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@                ���-��@��
�pV@        ��/����?
����M@        ��/����?H�4H�48@                H�4H�48@        ��/����?                ��/����?                ��/����?                        dJ�dJ�A@        0����/@�A�A>@        �cp>@                ��/����?�A�A>@                k�6k�69@        ��/����?��+��+@        ��/����?                        ��+��+@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��.hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhMh�hhK ��h��R�(KM��h��BH;         �                 �ꨣ?|��T�P�?-      5'�}@       �                 �<�?`1��>�?�       ���E�r@                          ҏ�?�4�����?�       �c_�Zr@                        �kΏ?�C P�}�?!       
YP.�J@                        �i?>">k�?       n�����D@                        ��%~?�k�G	�?       1@�8�C@                        �,=?�`@s'��?       ͡��[�@@       	                  h��?���3�?       ���(+�%@������������������������       �               �cp>@
                         l�@?���/��?       U��7�@                        `F|[?�d�$���?       �T�f@������������������������       �               ��/����?                        ��Km?      �<       ��#��@������������������������       �               ��#�� @������������������������       �               ��#�� @������������������������       �               �cp>@                        q�0?�B�� �?       �HI�7@                       ��z�?�(���?       x��uk!@������������������������       �               ��#���?������������������������       �      ��       ��/���@������������������������       �      ��	       ��|��,@                        ��!5?���/��?       @z$S��@������������������������       �               �cp>@������������������������       �               z�5��@                        �}?&�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?                        �u�?�Z�	7�?       j~���$@������������������������       �      �<       z�5��@������������������������       �      ��       ��/���@       �                 ��j�?��0+�'�?�       ��r�4n@        y                  ����?ʋ�r���?�       ���Y��l@!       `                 � �8?\��Y~
�?T       Ͽ����`@"       #                 0(\?��|G$�?:       ���=y�W@������������������������       �               ��b:��*@$       5                  �_�?$Sc�k�?3       �[Q�G(T@%       0                 �P�?{���[%�?       �I����8@&       -                 0��?^��jʄ�?
       @��m�0@'       ,                  P�"�?�m:�4�?       ���-X)@(       )                 @Ws�?��b�}�?       ���\�@������������������������       �               ��#�� @*       +                 x)�z?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �      ��       ��/���@.       /                  ���?�J���?       ��*]Y@������������������������       �               0#0# @������������������������       �               ��#�� @1       2                 �5�	? ����?       ��X�)B @������������������������       �               ��/����?3       4                 �{��?l����?       Q	K��@������������������������       �      �<       z�5��@������������������������       �      ȼ       ��/����?6       ]                 ��*?��>R��?$       �P��K@7       B                  ��&?(��ʀ�?!       r��I@8       A                    �?�PJo�x�?       T|qt�&@9       @                 �#h?����?       ��X�)B @:       ?                 ���>l����?       P	K��@;       >                 ;*��?����?       ��X�)B@<       =                F0qs?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �               z�5��@������������������������       �      ȼ       ��/����?������������������������       �      �<       �cp>@C       Z                 p]��?�"?���?       ���rD@D       S                  ᷁?�lMs���?       7�%}C@E       P                 �[�Z?�~�Hs=�?       ��?Z[0@F       O                 �U���p�T���?       ��e[�& @G       N                 �\��?JH����?       ��ϭ
*@H       M                 ��|?��Z�	7�?       j~���@I       L                 ��j�?�����?       ��X�)B@J       K                 `�sk?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?������������������������       �               0#0# @������������������������       �               ��#���?Q       R                  �Ab?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ���>��@T       U                 $^,W?����X��?       &��֞6@������������������������       �               ��/����?V       Y                 'uk?0 ����?       0
C>�5@W       X                 ��q�?��6L�n�?       �E#��h @������������������������       �      �<       ���>��@������������������������       �      ȼ       ��/����?������������������������       �      Լ       ��b:��*@[       \                 @�?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?^       _                 ����?      �<       ��/���@������������������������       �               ��/����?������������������������       �               �cp>@a       h                 0��?n��/��?       Г��OD@b       e                 p��?z�BG_��?       ���M�U3@c       d                 hf��>      �<       �cp>'@������������������������       �               ��/����?������������������������       �               /����/#@f       g                 �$9�?�ǧ\�?       �,W J@������������������������       �               H�4H�4@������������������������       �               0����/@i       p                 ��	�?��V�;�?       �(�A��4@j       k                  �_�?R�ђ���?       �oFݜh%@������������������������       �               0����/@l       m                  {X%?d%@�"�?       ��[�@������������������������       �               ��#���?n       o                 �+u?& k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      ��       ��/���@q       r                 ����?P-6���?       F��S=$@������������������������       �               ��#��@s       t                 �gY�?������?       ���'��@������������������������       �               0#0# @u       x                 � �?D��NV=�?       �t�ܲ@v       w                 `?��?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �      �<       ��/����?z       �                 Ў�?�TZf��?:       ��_�Y�W@{       �                  �?�
O�:��?        ��<�O�J@|       �                 ���r?��ș0��?       �6m�1zC@}       �                 �xK�?H�:V��?       �GP�A@~       �                 �y����	�� ��?       A�x��>@       �                 ���m?�����?       ��X�)B@�       �                   ��?bn����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �               ��b:��:@�       �                  pjS�?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@�       �                �3�q?�fm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?�       �                 P0Ы?4=�%�?
       t=�x�-@�       �                 ��Ղ?*µ*A
�?	       ��A抌)@�       �                 �-�?�(���?       y��uk!@�       �                 ��zk?      �<       ���-��@������������������������       �               ��/����?������������������������       �               �cp>@�       �                  �E�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                  ���?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@������������������������       �               ��#�� @�       �                 ?��? O�!]�?       ^��-c^D@�       �                 �30b?�w��d��?       �0���s+@�       �                 @1eQ? �Ϟi�?       ��ؠ�!@������������������������       �               ��/���@������������������������       �               ��+��+@�       �                 @Ax?���mf�?       毠�?b@������������������������       �      �<       ��/���@������������������������       �               0#0#�?�       �                 `<U�?����@��?       ;N,�;@�       �                 @X�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 pD�?r�cT�?       - w�8@�       �                 P��?r����?       Qz�i0@������������������������       �      ��	       ��8��8*@�       �                 p���?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 @��?T�4X��?       �<�?p�@�       �                 �*��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 t��I?Hy��]0�?       ���y"@�       �                 @-�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               0#0#@�       �                 ��?0�~:��?       �����)@������������������������       �               �C=�C=@�       �                 0"�?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �               0����/@�       �                 �1��?�*�'=P�?        �2"@������������������������       �               ��+��+@�       �                 �8��?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                 P� �?�}[W�R�?r       CB�+e@�       �                  (w�?�V&��o�?6       �Mj�R@�       �                 ��'s?"+(�UW�?/       �B~X"P@�       �                 ��N�?�+�b��?        �P��F@�       �                 <�Q?��l�?       ��.F�<@�       �                   ���?��$��?       @�"6@������������������������       �               �cp>@�       �                 0�,�?r��䭢�?       ^�[23@������������������������       �               ;��,��@�       �                  �E7?X�ih�<�?       ��
,@������������������������       �               vb'vb'"@�       �                 @���?hutee�?       Q9��@�       �                 �x�N?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �               0#0# @�       �                 p��U?��n��?       �-H�\@������������������������       �               ��/���@�       �                ༯U�?��q�R�?       C}Ԥ@������������������������       �               ��#���?�       �                 @6��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 �jU?��s`���?
       ���1�u0@�       �                 �C)�?Ǯ^���?       �.g���,@������������������������       �               0#0#�?������������������������       �               ��b:��*@�       �                ��1�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                  �"�?     ��<       ��)��)3@������������������������       �               0#0#�?������������������������       �               vb'vb'2@�       �                 ��N�?��XnP��?       ЭS`oM%@������������������������       �               ���-��@�       �                 P�*�?r�G���?       ��%�|@������������������������       �               ��/����?�       �                 �.K�?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�                        (��?��D�F�?<       ;�7���W@�       �                    �?D�T;���?#       >���hoJ@�       �                 ��A�?��"��?       <�x�LA@�       �                  -��?
�N���?       �3�R�E?@�       �                 �ƒ�?P-l�Fb�?       vrgN�3=@�       �                 `��?`.&��&�?       ��_B><@�       �                 ���?�����?       ��ȋ_)"@�       �                @u�/�?Hy��]0�?       ���y"@������������������������       �               ��/����?������������������������       �               ��+��+@�       �                 ���?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?������������������������       �        
       ��)��)3@������������������������       �      �<       ��/����?������������������������       �      ܼ       ��#�� @�       �                 @V�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?�                       \��?\G@^���?       X;�8�2@�       �                 ��?,�Z�K��?       X��Q�+@�       �                ��G�?�@G���?       hu��@������������������������       �               0#0#�?�       �                  �!�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?�                        ��=�?�@����?       ���a�#@������������������������       �               ��+��+@                      ���?hutee�?       Q9��@������������������������       �               ��/����?������������������������       �               H�4H�4@                       �w�?���mf�?       寠�?b@������������������������       �               �cp>@                       �r�?v�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?	                        s��?��Y�;�?       8�س��D@
                       �g<�?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?                      0��?      �<       vb'vb'B@������������������������       �               0#0#�?������������������������       �               dJ�dJ�A@�t�bh�hhK ��h��R�(KMKK��h �Bh  U^Cyc@.����/c@� � �d@Jy�5�_@u�����]@�+��+�K@Ky�5�_@�_��e�]@:k�6k�G@�P^Cy/@����z�A@0#0#�?�k(��"@�]�ڕ�?@0#0#�?��#�� @�]�ڕ�?@        ;��,��@��|��<@        ��#��@���-��@                �cp>@        ��#��@��/���@        ��#��@��/����?                ��/����?        ��#��@                ��#�� @                ��#�� @                        �cp>@        ��#���?h
��6@        ��#���?��/���@        ��#���?                        ��/���@                ��|��,@        z�5��@�cp>@                �cp>@        z�5��@                ��#���?        0#0#�?��#���?                                0#0#�?z�5��@��/���@        z�5��@                        ��/���@        .�����[@^�ڕ��T@(S2%S2G@.�����[@������S@��)��)C@��,���Q@e#6�aJ@#0#0&@$�}��O@�cp>�9@��+��+@��b:��*@                ~�5��H@�cp>�9@��+��+@;��,��$@�cp>'@H�4H�4@��#��@0����/#@H�4H�4@��#�� @0����/#@0#0#�?��#�� @��/����?0#0#�?��#�� @                        ��/����?0#0#�?                0#0#�?        ��/����?                ��/���@        ��#�� @        0#0# @                0#0# @��#�� @                z�5��@��/����?                ��/����?        z�5��@��/����?        z�5��@                        ��/����?        ������C@��|��,@0#0# @������C@鰑%@0#0# @z�5��@0����/@        z�5��@��/����?        z�5��@��/����?        z�5��@��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#�� @                z�5��@                        ��/����?                �cp>@        ��#��@@�cp>@0#0# @��#��@@��/���@0#0# @z�5��(@��/����?0#0# @��#��@��/����?0#0# @z�5��@��/����?0#0# @z�5��@��/����?        z�5��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                        ��/����?                        0#0# @��#���?                ��#�� @                ��#���?                ���>��@                <��,��4@��/����?                ��/����?        <��,��4@��/����?        ���>��@��/����?        ���>��@                        ��/����?        ��b:��*@                        ��/����?                ��/����?                ��/����?                ��/���@                ��/����?                �cp>@        ���>��@���-��:@H�4H�4@        On��O0@H�4H�4@        �cp>'@                ��/����?                /����/#@                0����/@H�4H�4@                H�4H�4@        0����/@        ���>��@鰑%@H�4H�4@��#�� @D�JԮD!@                0����/@        ��#�� @��/���@        ��#���?                ��#���?��/���@        ��#���?                        ��/���@        ;��,��@��/����?H�4H�4@��#��@                ��#���?��/����?H�4H�4@                0#0# @��#���?��/����?0#0#�?��#���?        0#0#�?                0#0#�?��#���?                        ��/����?        >��,��D@�cp>�9@�;�;;@��k(/D@���-��*@        Ey�5A@0����/@        ��#��@@��/����?        Kp�}>@��/����?        z�5��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ��#���?                ��b:��:@                z�5��@��/����?                ��/����?        z�5��@                ��#���?�cp>@                �cp>@        ��#���?                z�5��@D�JԮD!@        ��#��@D�JԮD!@        ��#���?��/���@                ���-��@                ��/����?                �cp>@        ��#���?��/����?                ��/����?        ��#���?                z�5��@��/����?                ��/����?        z�5��@                ��#�� @                ��#���?��On�(@�;�;;@        ��/���@H�4H�4@        ��/���@��+��+@        ��/���@                        ��+��+@        ��/���@0#0#�?        ��/���@                        0#0#�?��#���?0����/@��-��-5@        ��/����?0#0#�?                0#0#�?        ��/����?        ��#���?�cp>@��+��+4@        ��/����?�A�A.@                ��8��8*@        ��/����?0#0# @        ��/����?                        0#0# @��#���?��/����?��+��+@��#���?��/����?                ��/����?        ��#���?                        ��/����?��+��+@        ��/����?0#0#�?        ��/����?                        0#0#�?                0#0#@        0����/@0#0# @                �C=�C=@        0����/@0#0#�?                0#0#�?        0����/@                ��/����?0#0# @                ��+��+@        ��/����?H�4H�4@        ��/����?                        H�4H�4@z�5��8@�-����@@�+��+�[@<��,��4@0����/3@eJ�dJ�A@:��,��4@鰑%@B�A�@@<��,��4@鰑%@�C=�C=,@z�5��@/����/#@��8��8*@;��,��@0����/@H�4H�4(@        �cp>@        ;��,��@��/����?H�4H�4(@;��,��@                        ��/����?H�4H�4(@                vb'vb'"@        ��/����?H�4H�4@        ��/����?0#0#�?        ��/����?                        0#0#�?                0#0# @��#���?0����/@0#0#�?        ��/���@        ��#���?��/����?0#0#�?��#���?                        ��/����?0#0#�?        ��/����?                        0#0#�?���>��,@��/����?0#0#�?��b:��*@        0#0#�?                0#0#�?��b:��*@                ��#���?��/����?                ��/����?        ��#���?                                ��)��)3@                0#0#�?                vb'vb'2@        E�JԮD!@0#0# @        ���-��@                ��/����?0#0# @        ��/����?                ��/����?0#0# @        ��/����?                        0#0# @��#��@��|��,@�i��R@��#��@���-��*@fJ�dJ�A@��#��@0����/@k�6k�69@��#��@��/����?k�6k�69@��#�� @��/����?k�6k�69@��#�� @��/����?k�6k�69@��#�� @��/����?H�4H�4@        ��/����?��+��+@        ��/����?                        ��+��+@��#�� @        0#0#�?��#�� @                                0#0#�?                ��)��)3@        ��/����?        ��#�� @                        �cp>@                ��/����?                ��/����?                D�JԮD!@��+��+$@        0����/@vb'vb'"@        �cp>@0#0#�?                0#0#�?        �cp>@                ��/����?                ��/����?                ��/����?0#0# @                ��+��+@        ��/����?H�4H�4@        ��/����?                        H�4H�4@        ��/���@0#0#�?        �cp>@                ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?��+��+D@        ��/����?0#0#@                0#0#@        ��/����?                        vb'vb'B@                0#0#�?                dJ�dJ�A@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��~hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK݅�h��BX0         �                 ��\�?�-$��T�?       ��\�6}}@       y                   p��?$%y}�?�       �	�'�p@       <                 �vs?ق.t�?�       ��v�h3n@       )                 P^N<?JǱgw}�?I       ���c`@       "                  y��?�OH�V�?8       ��<+�Y@                        �U���fhK�4�?2       B�cp�W@                        �;�b?����a�?       �p�_��H@                        �c:?ذD���?	       ������6@	       
                 P���>)���?       y��uk!@������������������������       �               0����/@                        =�� ?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@                        `�u�?�_�A�?       肵�e`,@                         �Ur?���/��?       V��7�@������������������������       �               ��/����?                        �3�_?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �               z�5��@                           �?�(߫$��?       2H����:@                        ��s?X ����?       1
C>�5@������������������������       �               ��b:��*@                        @��x?��6L�n�?       �E#��h @������������������������       �               ��/����?������������������������       �      �<       ���>��@                         ��? 4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @                        �2�e?�q
<`&�?       ���g�F@������������������������       �               >��,��D@        !                 �X[Z?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@#       (                    �?�`���6�?       /u��֝!@$       '                 H�ӫ?���`�?       ��
�Me@%       &                 h�լ?r@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@������������������������       �               0#0# @������������������������       �               ��/����?*       ;                 �@	�?@�����?       ;-�s�V;@+       .                  `��?��\���?       �̑-`R9@,       -                 �Vp?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @/       :                 е�?�*d�^��?       ߌ�9�J6@0       3                 ��,b?�^�#΀�?       N�{��A5@1       2                 `n?f%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?4       9                  ��?�O
�*Q�?
       �͉V�M2@5       8                  ���?ʔfm���?       ��Z�N@6       7                 �ڡS?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      �<       ��|��,@������������������������       �      �<       ��#���?������������������������       �               0#0# @=       R                 �b�?�P���?J       h
���[@>       Q                  `<��?���SL:�?       5�.2�H@?       H                 �6O�?���#��?       �W�>H@@       G                 �x�.?��&���?       ��G2��<@A       F                 x��0?�`@s'��?
       Di_y,*+@B       E                 �p}?`n����?       � ��w<@C       D                 @��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#���?������������������������       �      ��       鰑%@������������������������       �               ��/���.@I       P                 ���? 6ׂ��?       �s�{ӎ3@J       O                 ��?�4�fP�?
       V���-@K       L                 �Ul?��q�R�?       C}Ԥ@������������������������       �               ��#���?M       N                 ��S�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               �cp>'@������������������������       �               ��+��+@������������������������       �      �<       ��#���?S       v                 �ju?�,��[�?+       �
��zN@T       q                 `��?.�LB��?%        b]��J@U       p                 5��?��,LP��?!       ��5�F@V       k                 pݔ�?��GӲ��?       �����B@W       d                 ��C?,)����?       <��3y�<@X       c                 ��U�? �e�>�?       n�B��3@Y       Z                ��'��?L[�Jg�?
       W�S0f�*@������������������������       �               ��/����?[       `                 �;�?��oR��?	       m�Q6�(@\       _                 �吂?P�k����?       a*pn�$@]       ^                 `��?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               ��#�� @a       b                 ���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               �cp>@e       j                 �΂�?: k�Lj�?       �q��l}#@f       i                 P:�?�(���?       y��uk!@g       h                 ����?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       ���-��@������������������������       �      �<       ��#���?l       o                 �-�;?R���'0�?       �C�� T"@m       n                 PL�?��6L�n�?       �E#��h @������������������������       �      �<       ���>��@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?������������������������       �               ���>��@r       u                 ���?�(���?       y��uk!@s       t                 �ڡC?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ���-��@w       x                    �?     ��<       �C=�C=@������������������������       �               H�4H�4@������������������������       �               0#0#@z       �                 Б�d?*��Ac�?       +t��-@{       ~                 ��j?���#��?       Z�f���'@|       }                   ���?|�r{��?       e�6� @������������������������       �               ���-��@������������������������       �               ��#���?       �                    �?�J���?       ��*]Y@������������������������       �               ��#�� @������������������������       �               0#0# @������������������������       �               H�4H�4@�       �                   s��?B.ܧ���?�       R1c�j@�       �                 P�|�?��']�?        7)� [H@�       �                     �?��c`�?       $��t5)@������������������������       �      ȼ       D�JԮD!@�       �                  �\�?̔fm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@�       �                 0�E�?�"�Hm��?       ,�N�B@�       �                 Ш��?��=����?       ~�(��p<@�       �                 ���?X�ih�<�?       ��
@������������������������       �               0#0#@�       �                 p
��?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 �nr�?(�b���?       �5��n5@�       �                 ����?���/��?       @z$S��@������������������������       �               z�5��@������������������������       �               �cp>@�       �                 `TF�?B� P?)�?       L.���.@�       �                   .p�?,Lj����?       ���T�,@������������������������       �               ���>��@�       �                 pq+�?��h��?       S�D'�@�       �                 `���?�J���?       ��*]Y@������������������������       �               ��#���?�       �                 ���?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               z�5��@������������������������       �               0#0#�?�       �                8���?�LU���?       i�ҹ^�@�       �                 �/�?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?������������������������       �               0����/@�       �                 pb\�?@$Ʉ|Z�?e       J�0��d@�       �                 `��\?,�����?U       �+��a@�       �                 �I��?|)vao��?/       ~�x�R@�       �                 NK�X?����K�?"       �f���K@�       �                   �0�?~�O<V��?       �S����6@�       �                 H��?Hy��]0�?       ���y"@������������������������       �               ��+��+@������������������������       �      ȼ       ��/����?�       �                 ��%�?������?
       3�<��0@�       �                  ����?<�a
=�?       ��l��+@������������������������       �               �cp>'@������������������������       �               0#0# @������������������������       �               H�4H�4@�       �                 @� ?4�z8o7�?       ,:����@@�       �                 �p�?\����?
       P	K��,@�       �                 JXˣ?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                  `���?pb8�Y�?       FJͰ(@������������������������       �      ��       ;��,��$@�       �                    �?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                  u�?A+2���?       ��1)3@�       �                 �н?D��15�?
       ��Qv�-@�       �                 �Ϻ�?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@�       �                 ��7�?�{����?       ـ�n�&&@������������������������       �               z�5��@�       �                 0���?����|e�?       �z �B�@�       �                  'T?`�ih�<�?       ��
@������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?������������������������       �               ��#��@�       �                 ����??�	,�?       >0�1b3@������������������������       �               ��/����?������������������������       �               S2%S2%1@�       �                 ����?0yAK;�?&       h�E�ׯN@�       �                 ����?0|�; -�?       ]��־�E@������������������������       �               ������C@�       �                    �?����|e�?       �z �B�@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?�       �                 ���?�*�'=P�?        �22@������������������������       �      �<       H�4H�4(@�       �                 ��k�?���`p��?       �����@������������������������       �               ��/����?������������������������       �      ��       0#0#@�       �                 �M�?`�v}�?       ���5>@�       �                 ��?X�ih�<�?       ��
@������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?�       �                    �?      �<       %S2%S27@������������������������       �               0#0# @������������������������       �               �A�A.@�t�bh�hhK ��h��R�(KK�KK��h �B�  ��b:��c@G:l��d@��jc@Np�}^@M!�M\@%S2%S27@�Gp�=]@��18�Z@vb'vb'2@���#8U@鰑E@0#0#@�b:���S@h
��6@0#0# @������S@On��O0@        Dy�5A@��/���.@        ZLg1��&@�cp>'@        ��#���?��/���@                0����/@        ��#���?�cp>@        ��#���?                        �cp>@        ;��,��$@��/���@        ��#��@��/���@                ��/����?        ��#��@��/����?                ��/����?        ��#��@                z�5��@                \Lg1��6@��/���@        ;��,��4@��/����?        ��b:��*@                ���>��@��/����?                ��/����?        ���>��@                ��#�� @�cp>@                �cp>@        ��#�� @                �GpAF@��/����?        >��,��D@                z�5��@��/����?                ��/����?        z�5��@                ��#���?�cp>@0#0# @��#���?0����/@0#0# @��#���?0����/@        ��#���?                        0����/@                        0#0# @        ��/����?        ;��,��@%jW�v%4@0#0# @;��,��@&jW�v%4@        ��#�� @��/����?                ��/����?        ��#�� @                z�5��@0����/3@        ��#�� @/����/3@        ��#���?��/����?                ��/����?        ��#���?                ��#���?D�JԮD1@        ��#���?�cp>@                �cp>@                ��/����?                ��/����?        ��#���?                        ��|��,@        ��#���?                                0#0# @���b:@@��P@�C=�C=,@��#��@������C@H�4H�4@z�5��@������C@H�4H�4@��#�� @���-��:@        ��#�� @�cp>'@        ��#�� @��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#���?                        鰑%@                ��/���.@        ��#���?��On�(@H�4H�4@��#���?��On�(@0#0#�?��#���?��/����?0#0#�?��#���?                        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>'@                        ��+��+@��#���?                ,�����;@��On�8@0#0# @,�����;@��On�8@0#0#�?��b:��:@E�JԮD1@0#0#�?������3@E�JԮD1@0#0#�?z�5��(@��/���.@0#0#�?<��,��$@��/���@0#0#�?<��,��$@��/����?0#0#�?        ��/����?        ;��,��$@��/����?0#0#�?�k(��"@        0#0#�?��#���?        0#0#�?                0#0#�?��#���?                ��#�� @                ��#���?��/����?                ��/����?        ��#���?                        �cp>@        ��#�� @��/���@        ��#���?��/���@        ��#���?��/����?                ��/����?        ��#���?                        ���-��@        ��#���?                ���>��@��/����?        ���>��@��/����?        ���>��@                        ��/����?                ��/����?        ���>��@                ��#���?��/���@        ��#���?��/����?                ��/����?        ��#���?                        ���-��@                        �C=�C=@                H�4H�4@                0#0#@z�5��@���-��@��+��+@z�5��@���-��@0#0# @��#���?���-��@                ���-��@        ��#���?                ��#�� @        0#0# @��#�� @                                0#0# @                H�4H�4@�YLg1B@��h
�G@?�C=ԃ`@��#��0@h
��6@��+��+$@��#���?�cp>'@                D�JԮD!@        ��#���?�cp>@        ��#���?                        �cp>@        �P^Cy/@鰑%@��+��+$@�P^Cy/@��/���@vb'vb'"@        ��/����?H�4H�4@                0#0#@        ��/����?0#0# @        ��/����?                        0#0# @�P^Cy/@�cp>@H�4H�4@z�5��@�cp>@        z�5��@                        �cp>@        z�5��(@        H�4H�4@z�5��(@        0#0# @���>��@                ;��,��@        0#0# @��#�� @        0#0# @��#���?                ��#���?        0#0# @��#���?                                0#0# @z�5��@                                0#0#�?        ���-��@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        0����/@        ������3@��On�8@*0#0�^@������3@�e�_��7@+S2%S2W@������3@鰑5@S2%S2%A@������3@0����/3@S2%S2%1@        ��On�(@��+��+$@        ��/����?��+��+@                ��+��+@        ��/����?                �cp>'@��+��+@        �cp>'@0#0# @        �cp>'@                        0#0# @                H�4H�4@������3@���-��@�C=�C=@z�5��(@��/����?        ��#���?��/����?        ��#���?                        ��/����?        \Lg1��&@��/����?        ;��,��$@                ��#���?��/����?                ��/����?        ��#���?                ���>��@0����/@�C=�C=@z�5��@0����/@�C=�C=@        �cp>@0#0#�?                0#0#�?        �cp>@        z�5��@��/����?H�4H�4@z�5��@                        ��/����?H�4H�4@        ��/����?H�4H�4@                H�4H�4@        ��/����?                ��/����?        ��#��@                        ��/����?S2%S2%1@        ��/����?                        S2%S2%1@        �cp>@�s?�s?M@        ��/����?��-��-E@                ������C@        ��/����?H�4H�4@                H�4H�4@        ��/����?                ��/����?0#0#0@                H�4H�4(@        ��/����?0#0#@        ��/����?                        0#0#@        ��/����?�s?�s?=@        ��/����?H�4H�4@                H�4H�4@        ��/����?                        %S2%S27@                0#0# @                �A�A.@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��.hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKՅ�h��B�.         �                 @E��? ud��O�?(      ��o��|}@       �                  �Mm�?ၟ;s�?�       ��Uk��t@       �                 0VҼ?tO$���?�       ���Cr@       w                 @��?�n����?�       mwF ��p@       t                  ���?������?�       j�{){l@       a                 0��?����"��?�       >�=�(j@       `                 `T��?��b��?o       lw�
ue@       ;                 �L�3?���#��?n       _1V�8e@	       :                 ��?�|̽R6�?A       � �I�Y@
       9                 pD	�?���F�Q�?=       ���%`/X@       0                 `JH~?�ۥܶ��?;       o�%2.wW@                        �l? ]A����?.       (>�-CS@                        �QZ?P�];�?       ��t�HA@                        ��aӾnzw��?       �B޳�X9@                        ��U?`n����?
       ����45@                        P���>���/��?       J9U6�+@������������������������       �               0����/@                        h�K?@���'0�?       �C�� T"@                        �$I�?|�6L�n�?       �E#��h @                          �x�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               z�5��@������������������������       �      ȼ       ��/����?������������������������       �      ��       ���>��@������������������������       �               ��#��@                         �"�?)���?       y��uk!@������������������������       �               ��#���?������������������������       �      �<       ��/���@       )                    �?�����_�?       ���FE@       (                 p'v�?�x�<�?       X&b��qA@        '                  ��q?���cE��?       b�co5@!       &                 �+"�?�3��F��?       mf9t{y4@"       #                 @�0�?�hK)�?       �h��K�2@������������������������       �               |�5��(@$       %                 �!�?�����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?������������������������       �      �<       ��/����?������������������������       �               ��b:��*@*       /                   \��?~��x���?       �!��4 @+       ,                 � �?D��NV=�?       �t�ܲ@������������������������       �               0#0#�?-       .                h�??f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#��@1       4                  �P��?��Sf\�?       i���0@2       3                 p���?�_�A�?       肵�e`@������������������������       �      �<       ;��,��@������������������������       �      ȼ       ��/����?5       8                 �؉�?\%��̫�?       �@�o#@6       7                 0d��?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               ��/���@������������������������       �      �       �cp>@������������������������       �               ���>��@<       W                 �<|�?_�̣�?-       b�X)P@=       @                  `��?hQ��?"       ��Я[[J@>       ?                 0�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#��@A       J                 ���@?x@ȱ��?       pm���SG@B       G                 Ы�q?�0��b�?
       SVl��0@C       F                 0�?���/��?       V��7�@D       E                  ���?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �               �cp>@H       I                    �?�(���?       y��uk!@������������������������       �               ��/���@������������������������       �               ��#���?K       L                 ����? �u�N��?       ������=@������������������������       �               :l��F:2@M       V                 ��֟?Ɣfm���?
       �0��z'@N       U                 �2*�?^%@�"�?	       �6�E�!@O       T                 `9�`?���/��?       @z$S��@P       S                 Pc	�?�Z�	7�?       j~���@Q       R                 �[�?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �      м       ��/����?������������������������       �      ȼ       �cp>@������������������������       �      �<       �cp>@X       _                 �d?��n?�?       �ZhiX�'@Y       ^                 �FX?��íxq�?       %2��-�@Z       ]                 pM�D?���mf�?       寠�?b@[       \                �Y���?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       �cp>@������������������������       �               ��#���?������������������������       �               H�4H�4@������������������������       �      �       H�4H�4@b       e                  ��3�?��m�'�?       Y��m�B@c       d                  `S��?l��H��?       v�I�@������������������������       �               z�5��@������������������������       �      �<       ��/���@f       s                 xV�}?n%��)��?       ,�ڈ�>@g       n                 �SR�?��ߐ��?       �X�(�<@h       i                 ��?��� ��?       �^�� @������������������������       �               ��/����?j       k                 PeT�?�djH�E�?       ^�\m�n@������������������������       �               ��#��@l       m                  Ц6�?x�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?o       p                 ���? �#�Ѵ�?       �)�B�4@������������������������       �               �k(��2@q       r                   \��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               0#0# @u       v                 ��}?�wV����?	       Bi�i�2@������������������������       �               ��#��0@������������������������       �               0#0# @x       �                 p���?(}�VuQ�?       ��C���E@y       z                 `iY�?((�V��?       Q�6Nv�B@������������������������       �               ��/���.@{       �                 pt��?��k���?       F+զm76@|       }                  ���?��٤ݸ?       ��<5�84@������������������������       �        
       D�JԮD1@~                        �۶�?f%@�"�?       ��[�@������������������������       �               ��/����?�       �                 �۲?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 0G�@?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 @���?���WW�?       �j�S@������������������������       �               z�5��@�       �                 (�r�?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                   �P�?�!��}�?       Ŷge��4@�       �                 ��?l@ȱ��?       nm���S'@������������������������       �      ��       0����/#@������������������������       �               ��#�� @�       �                 PGu�?t*�'=P�?        �2"@������������������������       �               H�4H�4@�       �                �\�ѓ?z��`p��?       �����@������������������������       �               0#0#�?�       �                 0�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 �i�?�C�����?       �^ť��E@�       �                 A}?��v��?       np��}27@�       �                 �m�?M�����?       p����.@�       �                 ����>���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      ��       ZLg1��&@�       �                 (�i<?�ǧ\�?       �,W J@������������������������       �      ��       0����/@������������������������       �               H�4H�4@�       �                  �y�?����|e�?       �L���3@�       �                 �u��?Jy��]0�?       �N-ۙ2@������������������������       �               ��+��+$@�       �                 ��?�~�&��?       ?�]��@������������������������       �               0#0#@�       �                 �0Md?�@G���?       hu��@�       �                  0p��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      м       ��/����?�       �                 �n��?h�p^w>�?S       ��4�a@�       �                   E(�?&��R��?<       ��c�	X@�       �                 p��?N�I��?	       tN���5@������������������������       �               ���-��@�       �                 �v�?�&��{*�?       z�����,@������������������������       �               �k(��"@������������������������       �               ��+��+@�       �                 �٠�?*�h����?3       K�o0�R@�       �                   �0�?Ơ)G�|�?$       i<I*�H@�       �                 `F �?�n�]:��?       ڸ����2@�       �                 y֩?���`p��?	       �����'@�       �                 ���?���mf�?       毠�?b@������������������������       �               �cp>@�       �                 0��?~�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ȼ       �C=�C=@�       �                 ��~?��|��?       ���ĺw@�       �                 �S|�?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               �cp>@�       �                 �{��?��p�?       ����>?@�       �                    �?����"�?       C��v7<@�       �                 p���?x����?       p�[50@������������������������       �               0#0# @�       �                 ��?z^�(���?       � K�h @�       �                 耯�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ȼ       H�4H�4@������������������������       �        	       H�4H�4(@�       �                  ���?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               k�6k�69@�       �                  �!�?�?�z�?       ��B,D@�       �                 �K��?�D#���?       �B�j@������������������������       �               0#0#@������������������������       �               ��#�� @�       �                 `�1�?�5���?       ��P9�A@������������������������       �               B�A�@@������������������������       �      �<       ��/����?�t�bh�hhK ��h��R�(KK�KK��h �B�  ��k(/d@��-��bd@���~�gb@��Gp_b@����-�a@;�;�F@�5�װ`@,����m`@�;�;;@�,���n`@0��18^@��)��)3@&�}��_@鰑U@S2%S2%1@�>��n[@鰑U@�A�A.@>��,��T@0����/S@H�4H�4(@>��,��T@0����/S@vb'vb'"@j1��tVQ@Pn��O@@0#0# @�P^CyO@Pn��O@@0#0# @�P^CyO@�_��e�=@0#0# @,�����K@&jW�v%4@0#0#�?������3@��|��,@        �k(��2@���-��@        ���>��,@���-��@        ���>��@���-��@                0����/@        ���>��@��/����?        ���>��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        z�5��@                        ��/����?        ���>��@                ��#��@                ��#���?��/���@        ��#���?                        ��/���@        �YLg1B@�cp>@0#0#�?�P^Cy?@��/���@        ��,���1@��/���@        ��,���1@�cp>@        ��,���1@��/����?        |�5��(@                ;��,��@��/����?        ;��,��@                        ��/����?                ��/����?                ��/����?        ��b:��*@                ;��,��@��/����?0#0#�?��#���?��/����?0#0#�?                0#0#�?��#���?��/����?        ��#���?                        ��/����?        ��#��@                z�5��@0����/#@0#0#�?;��,��@��/����?        ;��,��@                        ��/����?        ��#���?��/���@0#0#�?��#���?        0#0#�?                0#0#�?��#���?                        ��/���@                �cp>@        ���>��@                ��b:��*@h
��F@�C=�C=@|�5��(@'jW�v%D@        ��#��@��/����?                ��/����?        ��#��@                ��#�� @1����/C@        ;��,��@�cp>'@        ��#��@��/���@        ��#��@��/����?                ��/����?        ��#��@                        �cp>@        ��#���?��/���@                ��/���@        ��#���?                z�5��@���-��:@                :l��F:2@        z�5��@D�JԮD!@        z�5��@�cp>@        z�5��@�cp>@        z�5��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                        ��/����?                �cp>@                �cp>@        ��#���?��/���@�C=�C=@��#���?��/���@0#0#�?        ��/���@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@        ��#���?                                H�4H�4@                H�4H�4@��b:��:@��/���@H�4H�4@z�5��@��/���@        z�5��@                        ��/���@        �,����7@��/���@H�4H�4@�,����7@��/���@0#0#�?��#��@�cp>@0#0#�?        ��/����?        ��#��@��/����?0#0#�?��#��@                        ��/����?0#0#�?                0#0#�?        ��/����?        ������3@��/����?        �k(��2@                ��#���?��/����?        ��#���?                        ��/����?                        0#0# @��#��0@        0#0# @��#��0@                                0#0# @;��,��@;l��F:B@0#0# @��#�� @����z�A@                ��/���.@        ��#�� @&jW�v%4@        ��#���?0����/3@                D�JԮD1@        ��#���?��/����?                ��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#���?��/����?        ��#���?                        ��/����?        z�5��@��/����?0#0# @z�5��@                        ��/����?0#0# @        ��/����?                        0#0# @��#�� @鰑%@0#0# @��#�� @0����/#@                0����/#@        ��#�� @                        ��/����?0#0# @                H�4H�4@        ��/����?0#0# @                0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?��b:��*@�cp>'@vb'vb'2@��b:��*@���-��@H�4H�4@��b:��*@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ZLg1��&@                        0����/@H�4H�4@        0����/@                        H�4H�4@        0����/@�A�A.@        �cp>@�A�A.@                ��+��+$@        �cp>@��+��+@                0#0#@        �cp>@0#0#�?        �cp>@                ��/����?                ��/����?                        0#0#�?        ��/����?        ���>��,@'jW�v%4@z?�s?wY@z�5��(@/����/3@2#0#P@�k(��"@���-��@��+��+@        ���-��@        �k(��"@        ��+��+@�k(��"@                                ��+��+@z�5��@��On�(@����M@z�5��@��On�(@S2%S2%A@��#�� @E�JԮD!@0#0# @        ��/���@0#0# @        ��/���@0#0#�?        �cp>@                ��/����?0#0#�?        ��/����?                        0#0#�?                �C=�C=@��#�� @0����/@        ��#�� @��/����?                ��/����?        ��#�� @                        �cp>@        ��#���?��/���@��8��8:@��#���?��/����?��8��8:@��#���?��/����?�C=�C=,@                0#0# @��#���?��/����?H�4H�4@��#���?��/����?        ��#���?                        ��/����?                        H�4H�4@                H�4H�4(@        �cp>@                ��/����?                ��/����?                        k�6k�69@��#�� @��/����?�z��z�B@��#�� @        0#0#@                0#0#@��#�� @                        ��/����?B�A�@@                B�A�@@        ��/����?        �t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�DhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKم�h��Bx/         �                  b?��|*kO�?.      �����}@       �                 0CK�?�.y8���?�       ,�-��u@       r                 ��??om�YI��?�       �,���r@       ;                    �?$����?�       H�;!�=l@       :                 ��v�?�^ ҳ�?P       �x1u܁`@       /                 �ʨ�?P�'��?N       l3���_@       *                  �F�?.�l��?G       eg-��]@       #                  ���?�ފH/3�?A       �$�zZ[@	                         L��?����,��?(       �{u;y�M@
                         `S��?���?       jz3��9@������������������������       �               ��/����?                          ��?�6�%�?       t��Ce�8@                        г��?@ ����?       1
C>�5@������������������������       �      ��	       ������3@                        ��aӾ���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?                        �/��?R����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?                        p|�o?�\�sF��?       W>��A@                        @I��>R�ђ���?       �oFݜh%@������������������������       �               ��/���@                             ��|��?       ���ĺw@                        Z�K?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               �cp>@                        @�u?΃�\��?       �D+զm7@������������������������       �               <��,��$@       "                �Su�z?��?	       ��l}�'*@        !                 ���?8�c3���?       �uk��!@������������������������       �               0����/@������������������������       �               ��#��@������������������������       �               ��#��@$       )                 P�ּ?X[�T��?       yԼ|�H@%       &                 `�?�M2�8ӣ?       h�R�dIH@������������������������       �               �k(���E@'       (                  �u��?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �      ��       0#0#�?+       ,                 ����?P��H��?       v�I�@������������������������       �               �cp>@-       .                   +Y�?����?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?0       5                  �t�?[n���2�?       HX-�[�%@1       4                 0�qw?�`@s'��?       Ei_y,*@2       3                @0W=e?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �               ��/���@6       7                  9e�?�zœ���?       IG���t@������������������������       �               ��#�� @8       9                 ��{�?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               0����/@<       =                  `<��?+<X���?;       l�X7xW@������������������������       �               0����/@>       K                 tlq?؎�6��?8       ���l9EV@?       F                 @���?��/ʪ��?	       H�Ų��1@@       C                 �m۶?,��c`�?       &��t5)@A       B                 �m�?$ k�Lj�?       �q��l}@������������������������       �               ��/���@������������������������       �      м       ��#���?D       E                 �!P?      �<       ��/���@������������������������       �               �cp>@������������������������       �               0����/@G       J                 .�X?�d�$���?       �T�f@H       I                 ��� ?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      ��       ��#�� @L       g                 �^Ҧ?���/u�?/       h;3@��Q@M       d                 `���?�X�@K�?"       g���luI@N       c                 �!�?��j�:��?       O�_E:@O       \                 �sf�?aTi�<��?       	���8@P       Q                 @��>�Z��.��?       .���d.@������������������������       �               ��/����?R       W                 `Ԙ�?�mh�y<�?       D��y,@S       V                 @�n�>�FO���?       �ߌ$@T       U                 �=��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ��       ��#�� @X       [                 P�L�?B��NV=�?       �t�ܲ@Y       Z                 �И�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               ��#���?]       b                ���[�?j%@�"�?       �6�E�!@^       _                  ���?ʔfm���?       ��Z�N@������������������������       �               ��#���?`       a                 �@�?�`@s'��?       Ei_y,*@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               0#0# @e       f                 �كv?      �<       |�5��8@������������������������       �               ��#���?������������������������       �               �,����7@h       m                 ��2�?:&��:��?       ��0kk�4@i       j                  �G?�?@W���?       �$!��.@������������������������       �               鰑%@k       l                 �~��?jutee�?       Q9��@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?n       o                 ��@�?@�N9���?       ��{j�@������������������������       �               ��#���?p       q                  �9��?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@s       �                 ��U�?uM�~L�?2       �1�j�R@t       �                  ����?���Z�)�?$       �d���K@u       x                  �X?ҿCB�?       �[�xA@v       w                 @�Ks?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@y       ~                 P�N�?&t���?       Ŷ���=@z       {                  �x��?�B�� �?       �HI�7@������������������������       �               D�JԮD1@|       }                 ���R?t@ȱ��?       om���S@������������������������       �               0����/@������������������������       �               ��#���?       �                 `}��?��r�g��?       ��1ֻ�@�       �                 �N��?T����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �               �cp>@�       �                 ��D�?�|���Y�?       �~��95@�       �                 �!�?z��`p��?       �����@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?�       �                 ���>�˝Ѝ��?	       b����.@������������������������       �               0#0#�?�       �                 p�D�?�B���?       F��,�,@�       �                 P��t?tb8�Y�?       FJͰ(@�       �                 ��dp?����?       ��X�)B@������������������������       �      ��       z�5��@������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?�       �                 p��?h[nD���?       ���y�O3@������������������������       �      ��       On��O0@�       �                    �?��q�R�?       C}Ԥ@������������������������       �               ��#���?�       �                 �^c�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 |�L?X7��{N�?$       �����fI@�       �                 P7J�?��w(�?       -�,?/>@�       �                 ����?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                    �?����"�?       C��v7<@�       �                 ���?1����?       �`O��"@������������������������       �               ��+��+@�       �                 ��?�3`���?       -�r��@�       �                 0�̱?��q�R�?       C}Ԥ@�       �                  w�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               0#0#�?�       �                  P���?      �<       ��)��)3@������������������������       �               0#0#�?������������������������       �        
       vb'vb'2@�       �                 �m��?��7�W��?       �S]��4@�       �                  ���? �Ϟi�?       
��ؠ�!@������������������������       �               ��/���@������������������������       �      ȼ       ��+��+@�       �                 p�A�?Δfm���?	       �0��z'@�       �                    �?�ۜ�x�?       d��إV#@������������������������       �               0����/@�       �                 y��?  k�Lj�?       �q��l}@������������������������       �      �<       ��/���@������������������������       �               ��#���?������������������������       �               ��#�� @�       �                 �ֈ?��Ց�?M       �>Z6K^@�       �                 @F�|�ҭ�x�?       �
�H��0@������������������������       �               �cp>@�       �                 �۶�?F�Uέ��?
       Bq��+@�       �                  2�z?�D�-,�?       �D'ŰO@�       �                 �E3[?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               H�4H�4@�       �                 �ܳ?z�G���?       ��%�|@������������������������       �               �cp>@�       �                 �8��?�@����?       ���a�@�       �                 �@�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       H�4H�4@�       �                 �j�}?|}/A{E�?A       V�( AZ@�       �                 ��p?nutee�?       �UY���-@������������������������       �               vb'vb'"@������������������������       �               �cp>@�       �                 �qҍ?�$^F��?:       ��]��`V@�       �                 pT��?�g���E�?       �m���9@�       �                 `�4x?�w��Z��?       �R9@�       �                 @�:�?�T`�[k�?	       �m����0@�       �                 �lw?��E�B��?       dߞKC.@�       �                  ���?t��ճC�?       y��l$,@������������������������       �               ��+��+$@�       �                   Y��?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?������������������������       �               0#0# @������������������������       �      �<       ��/����?�       �                 (���?      �<*       R��N��O@������������������������       �               0#0# @������������������������       �        )       /��+��N@�t�b��     h�hhK ��h��R�(KK�KK��h �BX  cCy��d@�[<���b@�؉��Ic@Qg1���d@����/�`@�˷|˷I@	��GPd@�_��e�]@��)��)3@������a@����z�Q@H�4H�4(@ZUUUU�X@��/���>@H�4H�4@ZUUUU�X@�cp>�9@H�4H�4@�t�Y�W@&jW�v%4@0#0# @^Lg1��V@On��O0@0#0# @�k(���E@��/���.@0#0#�?\Lg1��6@��/����?0#0#�?        ��/����?        \Lg1��6@��/����?0#0#�?<��,��4@��/����?        ������3@                ��#���?��/����?                ��/����?        ��#���?                ��#�� @        0#0#�?��#�� @                                0#0#�?>��,��4@���-��*@        ��#�� @D�JԮD!@                ��/���@        ��#�� @0����/@        ��#�� @��/����?        ��#�� @                        ��/����?                �cp>@        �k(��2@0����/@        <��,��$@                ��#�� @0����/@        ��#��@0����/@                0����/@        ��#��@                ��#��@                �,����G@��/����?0#0#�?�,����G@��/����?        �k(���E@                ��#��@��/����?        ��#��@                        ��/����?                        0#0#�?z�5��@��/���@                �cp>@        z�5��@��/����?        z�5��@                        ��/����?        ��#��@�cp>@0#0#�?��#���?�cp>@        ��#���?��/����?                ��/����?        ��#���?                        ��/���@        z�5��@        0#0#�?��#�� @                ��#���?        0#0#�?                0#0#�?��#���?                        0����/@        �GpAF@'jW�v%D@vb'vb'"@        0����/@        �GpAF@����z�A@vb'vb'"@;��,��@��On�(@        ��#���?�cp>'@        ��#���?��/���@                ��/���@        ��#���?                        ��/���@                �cp>@                0����/@        ��#��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ��#�� @                ������C@�cp>7@vb'vb'"@d:��,&C@0����/#@H�4H�4@��b:��*@0����/#@H�4H�4@��b:��*@0����/#@0#0#�?<��,��$@��/���@0#0#�?        ��/����?        <��,��$@�cp>@0#0#�?�k(��"@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                ��#���?��/����?0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?        ��#���?                z�5��@�cp>@        ��#�� @�cp>@        ��#���?                ��#���?�cp>@        ��#���?                        �cp>@        ��#���?                                0#0# @|�5��8@                ��#���?                �,����7@                ��#���?���-��*@H�4H�4@        ��On�(@H�4H�4@        鰑%@                ��/����?H�4H�4@                H�4H�4@        ��/����?        ��#���?��/����?H�4H�4@��#���?                        ��/����?H�4H�4@        ��/����?                        H�4H�4@������3@�e�_��G@�C=�C=@�k(��2@��/���>@H�4H�4@���>��@�cp>�9@0#0#�?��#��@��/����?                ��/����?        ��#��@                z�5��@��On�8@0#0#�?��#���?h
��6@                D�JԮD1@        ��#���?0����/@                0����/@        ��#���?                ��#�� @�cp>@0#0#�?��#�� @        0#0#�?                0#0#�?��#�� @                        �cp>@        [Lg1��&@0����/@��+��+@        ��/����?0#0#@                0#0#@        ��/����?        ZLg1��&@�cp>@0#0#�?                0#0#�?[Lg1��&@�cp>@        [Lg1��&@��/����?        z�5��@��/����?        z�5��@                        ��/����?        ��#�� @                        ��/����?        ��#���?E�JԮD1@0#0#�?        On��O0@        ��#���?��/����?0#0#�?��#���?                        ��/����?0#0#�?        ��/����?                        0#0#�?��#��@��|��,@0#0#@@��#���?��/����?�;�;;@        ��/����?0#0#�?                0#0#�?        ��/����?        ��#���?��/����?��8��8:@��#���?��/����?�C=�C=@                ��+��+@��#���?��/����?0#0# @��#���?��/����?0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?��#���?                                0#0#�?                ��)��)3@                0#0#�?                vb'vb'2@z�5��@��On�(@��+��+@        ��/���@��+��+@        ��/���@                        ��+��+@z�5��@E�JԮD!@        ��#���?E�JԮD!@                0����/@        ��#���?��/���@                ��/���@        ��#���?                ��#�� @                ��#���?E�JԮD1@�˷|˷Y@��#���?���-��@vb'vb'"@        �cp>@        ��#���?��/���@vb'vb'"@��#���?        ��+��+@��#���?        0#0# @��#���?                                0#0# @                H�4H�4@        ��/���@0#0#@        �cp>@                ��/����?0#0#@        ��/����?0#0#�?        ��/����?                        0#0#�?                H�4H�4@        鰑%@2��-�rW@        �cp>@vb'vb'"@                vb'vb'"@        �cp>@                0����/@��-��-U@        0����/@��-��-5@        ��/���@��-��-5@        ��/���@��8��8*@        ��/����?��8��8*@        ��/����?��8��8*@                ��+��+$@        ��/����?H�4H�4@        ��/����?                        H�4H�4@        ��/����?                ��/����?                        0#0# @        ��/����?                        R��N��O@                0#0# @                /��+��N@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ���MhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKυ�h��BH-         �                 ���b?P0�T�?)      C����}@       �                 �B��?p�2(��?�       �ۆ59�u@       \                 `��?�S�ߐ�?�       $����{p@       Q                 ��~?�p?2�?{       K�ƴ�6g@       B                 ���@?c�z��K�?i       ��E��c@       ;                 /O�?�K��_��?S       v��ZU_@       (                 �U���:2
����?L       �3?��M]@                        pe�S?(���R�?(       6�jAJ�L@	                        `:e?��\���?       �̑-`R9@
                        p���>�4��v�?
       �Y-"�'@                        .25Q?l@ȱ��?       nm���S@                        ��V?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ��       ��/���@                        �Z�?bn����?       � ��w<@                         8hV?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               ��#�� @                        P\�>      �<       ���-��*@������������������������       �               ��/����?������������������������       �               ��On�(@       %                 �3�_?���?       ���*@@                        �'�?
�kO���?       �y�ڲ�9@������������������������       �               z�5��@                        P�^�?����]L�?       O66�ͯ3@                         ��j?)���?       y��uk!@������������������������       �               ��#���?������������������������       �               ��/���@       $                    �?�ݛ��4�?       $�V�%�%@        #                   +Y�?C��X�&�?       �6��	�@!       "                   �0�?�zœ���?       IG���t@������������������������       �               z�5��@������������������������       �               0#0#�?������������������������       �      �<       ��/���@������������������������       �               H�4H�4@&       '                  ��? ����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?)       8                 �u�?�ө@h�?$       �����M@*       5                 1[v?��@����?!       ��`�L@+       4                 ���X?�I��X[�?       �h��G@,       -                 8Q�S?T�؈�w�?       q���S#G@������������������������       �               ��/����?.       3                 P��1?`�+(�s�?       �9Շ�F@/       0                 @��?��E�B��?       �'�xr�6@������������������������       �               �P^Cy/@1       2                 ��=�?�)z� ��?       �\�@������������������������       �               �cp>@������������������������       �               ��#��@������������������������       �               [Lg1��6@������������������������       �      �<       ��/����?6       7                 ��A�?vQ��?       �s�=�!@������������������������       �      ��       ���-��@������������������������       �               ��#�� @9       :                 p��1?      �<       ��/���@������������������������       �               ��/����?������������������������       �               �cp>@<       =                 �D��?�,���O�?       ���/> @������������������������       �               H�4H�4@>       A                  �p�?     ��?       "F�b@?       @                 j�1�?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?������������������������       �               0#0# @C       P                 �(i�?��f^�|�?       ��S�^u@@D       O                  .Dy?|�K�m��?       S�D]�>@E       H                 p��g? ���w��?       �"�!-�=@F       G                ��fr�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?I       J                  ���?��XG�J�?       m����;@������������������������       �               鰑5@K       L                 X?�`@s'��?       Ei_y,*@������������������������       �               ��/���@M       N                 ��f?d%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �               0#0# @R       W                 �l�?|	T��?        ��ew;@S       T                 ����?0 ����?       2
C>�5@������������������������       �               \Lg1��&@U       V                  �^�?�FO���?       �ߌ$@������������������������       �               ��/����?������������������������       �               �k(��"@X       Y                 ����?�֪u�_�?       ��?�8@������������������������       �               �cp>@Z       [                 P4��?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?]       ~                 pM�D?&h�c��?6       �q�hS�S@^       _                 ��r<?\9TNb��?.       ��ȥQ@������������������������       �               ��/����?`       u                  ��^�?У.�1�?-       MDJ�ٕP@a       p                 �&�?XL�Е��?$       ���*�K@b       c                 ���?�G|:=*�?        �`���G@������������������������       �               ��,���1@d       g                   ��?>i1�Z��?       ��g���=@e       f                 ����?2�c3���?       �uk��!@������������������������       �               0����/@������������������������       �               ��#��@h       o                 0�� ?Ț����?       �ڬ�ڬ4@i       n                  @?��? �%�?        ����.@j       m                  C�?�zœ���?       IG���t@k       l                pn�ǣ?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �      ��       [Lg1��&@������������������������       �               ;��,��@q       r                 �U�<?��V���?       �0��M @������������������������       �               ;��,��@s       t                 �{��?���`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @v       w                 ة q?E
:����?	       {��"�%@������������������������       �               ��#�� @x       }                  `<��?���1n�?       =���4�!@y       z                 �K�?�֪u�_�?       ��?�8@������������������������       �               ��/���@{       |                 �m��?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               z�5��@       �                 @� %?  k�Lj�?       �q��l}#@������������������������       �               ��#���?�       �                 �˱?)���?       y��uk!@������������������������       �               0����/@�       �                 �s%�?Ȕfm���?       ��Z�N@������������������������       �               ��#���?�       �                 Њ�H?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?�       �                 �Zz�?����d��?0       �����T@�       �                 x��?��%�f��?       TB�a�H@�       �                  1��?����|e�?       �z �B�@������������������������       �               ��+��+@�       �                 P�o�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 -��?���M��?       �2N	�D@�       �                 �Q��?F��3��?       �_q>c3@�       �                 px��?�0�~��?
       r��GQ1@������������������������       �        	       On��O0@������������������������       �               0#0#�?������������������������       �      �<       ��#�� @�       �                    �?�ن�f�?       Y+4�4@�       �                8�|�?r^�(���?       � K�h @�       �                 A��?P�ih�<�?       ��
@������������������������       �               0#0#@�       �                 ���?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               ��#���?�       �                  l�V?~-�E�T�?       ��<)@�       �                  s��?�}	;	�?       vK�>4%@������������������������       �               D�JԮD!@�       �                 �9/�?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               0#0# @�       �                 pw��?zn����?       ��ۥz�A@�       �                  ���?���)��?       U���*7@�       �                 @�ٲ?H��aB��?	       ����2@�       �                ����}?�`���6�?       /u��֝!@�       �                 �u�?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?�       �                 ��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               0����/@������������������������       �      ��       �k(��"@������������������������       �               ��+��+@�       �                �{\��?      �<       H�4H�4(@������������������������       �               vb'vb'"@������������������������       �               H�4H�4@�       �                 0�0�?�柞��?H       �إM_@�       �                 0#ή?��3A+B�?       ��ɪmE@�       �                 ��Wv?$�[tq�?       ��'�~)@�       �                  gm?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@�       �                 x�׀?�;[��G�?       �O�;�]!@������������������������       �      �<       ��/���@������������������������       �               0#0#�?�       �                 0٘�?�?�0�!�?       ��G�>@�       �                 @��?lutee�?       Q9��@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                 0��?�-�bƲ?       >�7*9@�       �                 ���?�^�F�M�?       ��ޚ�&@������������������������       �               ��+��+$@������������������������       �      ȼ       ��/����?�       �                 �zW�?      �<       �C=�C=,@������������������������       �               0#0# @������������������������       �               H�4H�4(@�       �                    �?hC-m#,�?1       ��EsЖT@������������������������       �               T2%S2%A@�       �                 @�-�?H
����?       *f�nH@������������������������       �      м       k�6k�69@�       �                  �j�?��9 ���?       �z��)�6@�       �                 �%{�?��^���?       ���w!@������������������������       �      ��       ���-��@������������������������       �               0#0# @������������������������       �               �C=�C=,@�t�bh�hhK ��h��R�(KK�KK��h �Bh  �>��d@	鰑Nc@������c@������c@��t�Ha@������J@�}��a@i��F:lY@vb'vb'2@:��P^�V@��-��bT@�C=�C=,@k1��tVQ@r�'�x�R@��8��8*@"�}��P@�e�_��G@��+��+$@�P^CyMP@�e�_��G@0#0#@<��,��4@Pn��O@@0#0#@;��,��@%jW�v%4@        ;��,��@���-��@        ��#���?0����/@        ��#���?��/����?        ��#���?                        ��/����?                ��/���@        ��#��@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ��#�� @                        ���-��*@                ��/����?                ��On�(@        �P^Cy/@��On�(@0#0#@<��,��$@�cp>'@0#0#@z�5��@                ��#��@�cp>'@0#0#@��#���?��/���@        ��#���?                        ��/���@        z�5��@��/���@0#0#@z�5��@��/���@0#0#�?z�5��@        0#0#�?z�5��@                                0#0#�?        ��/���@                        H�4H�4@;��,��@��/����?        ;��,��@                        ��/����?        �GpAF@��/���.@        �GpAF@�cp>'@        ���#8E@0����/@        ���#8E@��/���@                ��/����?        ���#8E@�cp>@        ������3@�cp>@        �P^Cy/@                ��#��@�cp>@                �cp>@        ��#��@                [Lg1��6@                        ��/����?        ��#�� @���-��@                ���-��@        ��#�� @                        ��/���@                ��/����?                �cp>@        ��#�� @        H�4H�4@                H�4H�4@��#�� @        H�4H�4@��#�� @        0#0#�?��#�� @                                0#0#�?                0#0# @��#�� @�a#6�;@H�4H�4@��#�� @�a#6�;@0#0#�?��#�� @�a#6�;@        ��#���?��/����?                ��/����?        ��#���?                ��#���?���-��:@                鰑5@        ��#���?�cp>@                ��/���@        ��#���?��/����?        ��#���?                        ��/����?                        0#0#�?                0#0# @<��,��4@�cp>@0#0#�?<��,��4@��/����?        \Lg1��&@                �k(��"@��/����?                ��/����?        �k(��"@                        0����/@0#0#�?        �cp>@                ��/����?0#0#�?        ��/����?                        0#0#�?��b:��J@%jW�v%4@0#0#@�#���I@��On�(@0#0#@        ��/����?        �#���I@鰑%@0#0#@����JG@�cp>@H�4H�4@>��,��D@0����/@0#0#�?��,���1@                �,����7@0����/@0#0#�?��#��@0����/@                0����/@        ��#��@                ������3@        0#0#�?���>��,@        0#0#�?z�5��@        0#0#�?��#���?        0#0#�?                0#0#�?��#���?                ��#�� @                [Lg1��&@                ;��,��@                ;��,��@��/����?0#0# @;��,��@                        ��/����?0#0# @        ��/����?                        0#0# @;��,��@0����/@0#0#�?��#�� @                z�5��@0����/@0#0#�?        0����/@0#0#�?        ��/���@                ��/����?0#0#�?        ��/����?                        0#0#�?z�5��@                ��#�� @��/���@        ��#���?                ��#���?��/���@                0����/@        ��#���?�cp>@        ��#���?                        �cp>@                ��/����?                ��/����?        ��b:��*@F�JԮDA@dJ�dJ�A@z�5��@��|��<@0#0#0@        ��/����?H�4H�4@                ��+��+@        ��/����?0#0#�?                0#0#�?        ��/����?        z�5��@���-��:@��+��+$@��#�� @On��O0@0#0#�?        On��O0@0#0#�?        On��O0@                        0#0#�?��#�� @                ��#���?鰑%@vb'vb'"@��#���?��/����?H�4H�4@        ��/����?H�4H�4@                0#0#@        ��/����?0#0# @        ��/����?                        0#0# @��#���?                        0����/#@H�4H�4@        0����/#@0#0#�?        D�JԮD!@                ��/����?0#0#�?        ��/����?                        0#0#�?                0#0# @;��,��$@�cp>@��)��)3@;��,��$@�cp>@�C=�C=@<��,��$@�cp>@0#0# @��#���?�cp>@0#0# @��#���?        0#0# @                0#0# @��#���?                        �cp>@                ��/����?                0����/@        �k(��"@                                ��+��+@                H�4H�4(@                vb'vb'"@                H�4H�4@z�5��@:l��F:2@�Wx�W�Y@z�5��@�cp>'@�C=�C=<@z�5��@D�JԮD!@0#0#�?z�5��@��/����?                ��/����?        z�5��@                        ��/���@0#0#�?        ��/���@                        0#0#�?        �cp>@�;�;;@        ��/����?H�4H�4@        ��/����?                        H�4H�4@        ��/����?H�4H�48@        ��/����?��+��+$@                ��+��+$@        ��/����?                        �C=�C=,@                0#0# @                H�4H�4(@        ���-��@�i��R@                T2%S2%A@        ���-��@�ڬ�ڬD@                k�6k�69@        ���-��@0#0#0@        ���-��@0#0# @        ���-��@                        0#0# @                �C=�C=,@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ9M�hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK߅�h��B�0         �                 pK�b?Z�Αx9�?      �7��Ɩ}@       �                 `m�?�N�0��?�        ��3�u@       �                 P7&E?�=Sbe��?�       cr"(��q@       a                 �U����= �?�       �>�ų�m@       L                  ����?��h�+?�?^       �CfA��a@       %                 ���?���?H       gZc��Z@                        P¤X?��A�7��?"       �2�mqF@                         �g<�?��/ʪ��?       H�Ų��1@	                         @��?�^�#΀�?       O�{��A%@
                         pjS�?      �<       0����/@������������������������       �               ��/����?������������������������       �               ��/���@                        0+��>r@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@                        �$I�?�)z� ��?       �\�@������������������������       �               ��#�� @                        @I��>
4=�%�?       �(J��@������������������������       �               ��/����?                        ���`?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @                         �.�?�����?       R�T3;=;@                        ��t?d�T��?       ��R�)@������������������������       �               ��#��@                          ҏ�?)���?       y��uk!@������������������������       �               0����/@                        p܀�?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@       $                 �~��?��DNpk�?       �k�Z$�,@        !                 𪛀?X�s�	�?       f���*@������������������������       �               z�5��@"       #                 �5��?L����?       P	K��@������������������������       �               ��/����?������������������������       �               z�5��@������������������������       �               0#0#�?&       =                   s��?�M����?&       ��Ӫ�N@'       (                  �ß?��4�,��?       /�i0�@@������������������������       �               0#0#@)       :                   \��?(�6N�?       ��ʲ�!=@*       /                 p���?\�����?       ��d�?K9@+       .                 [�?����]L�?       N66�ͯ@,       -                 h�լ?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               �cp>@0       1                  ��g�?�*A� f�?       fT�L_4@������������������������       �               ��/����?2       9                 `(��?�Ͳ�S{�?       pս��i3@3       8                  n��?�����?       N��o�g2@4       7                 0�0�?�����?       �Ä�>c(@5       6                  �P��?�FO���?       �ߌ$@������������������������       �               �k(��"@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?������������������������       �               z�5��@������������������������       �               0#0#�?;       <                 @�W�?      �<       ��/���@������������������������       �               ��/����?������������������������       �               �cp>@>       I                 �4�?n��UTH�?       �Yzh��<@?       H                 �Zx�?.�(��?       ��V-�:@@       A                 �~�?Н�/U��?       �+�f��9@������������������������       �               0#0# @B       G                 pI�?�q�Ptܳ?       P�� 5�7@C       D                   ��?X�j���?       ���z"@������������������������       �               z�5��@E       F                  ���?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      �<       ���>��,@������������������������       �      �<       ��/����?J       K                 ��?��G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?M       ^                  @�a�?�~���;�?       .��>8�A@N       S                 p'v�?F�Ӊa��?       U����3@@O       R                 `#z?e��}�?	       ��Se+@P       Q                    �?r@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@������������������������       �      �<       ��/���@T       U                 �p�?��X\��?       ��BM��2@������������������������       �               H�4H�4@V       [                  ���?�V�J��?       �Uk�T�)@W       Z                 ��i-?p�r{��?       e�6� @X       Y                    �?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               0����/@\       ]                ���u?    ��?       "F�b@������������������������       �               H�4H�4@������������������������       �               ��#�� @_       `                 ��'�?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ��#�� @b       {                 �~��?�8����?8       ��?zW@c       f                  ��>�x�<�?)       Z&b��qQ@d       e                ��l�~?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?g       z                 ����?X�4ƺ&�?'       ��%��P@h       m                 �kd1?l҃l[ �?%       ǻ���NN@i       j                 �x?��+�*�?       wȚ�
A@������������������������       �               �P^Cy?@k       l                  Pmj�?dn����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?n       o                 P��1?���&���?       ���[��:@������������������������       �               ��/����?p       u                 (6e?��6L�n�?       ��4}i�8@q       r                 �p�?�N:�*ط?       I�G�3@������������������������       �      ��       ���>��,@s       t                 88�s?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?v       w                  ��j?�Z�	7�?       j~���@������������������������       �               ��#�� @x       y                 Ȯ�?f%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �               z�5��@|                         �3?£���c�?       �>�!J!8@}       ~                 ����?��[����?       Hl�_A@������������������������       �               0����/@������������������������       �               0#0# @�       �                 0*tC?v�w�o�?       �c/�P1@������������������������       �               <��,��$@�       �                 �΂�?��R��?       y:b|�@�       �                 P4��?wT �+��?       ��>Y��@�       �                 �j{?Ȕfm���?       ��Z�N@������������������������       �               ��/����?�       �                 �:h�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               0#0# @������������������������       �               ��#���?�       �                 ��U�?���W�1�?       ��)��G@�       �                 �7�?�a�Q��?       ���nݔ?@�       �                 ��? ��c`�?       %��t5)@������������������������       �      ��       E�JԮD!@�       �                  p�Z?̔fm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@�       �                 ���>$�e�>�?       n�B��3@������������������������       �               0#0#�?�       �                 �~ɀ?� �_rK�?       J�@��2@�       �                    �?$ k�Lj�?       �q��l}@������������������������       �               ��/���@������������������������       �      м       ��#���?�       �                 ��8�?�3���r�?
       ��7�nN*@�       �                 0�H�?�)z� ��?       �\�@������������������������       �               ��/����?�       �                 ��I�?�d�$���?       �T�f@������������������������       �               z�5��@�       �                    �?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                  �h�?�����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?�       �                  `%+�?      �<	       Nn��O0@������������������������       �               �cp>@������������������������       �               ���-��*@�       �                 �%�?b<B�
��?&       ��{iBP@�       �                 H=	�?X�Z�E��?       ���H@�       �                 `��u?��N��?	       B5ٴ[Z0@������������������������       �               0#0#@�       �                 �X\�?��oR��?       l�Q6�(@�       �                 @eb�?l7Y���?       ���r�&@������������������������       �               0#0#�?������������������������       �               <��,��$@������������������������       �      ȼ       ��/����?�       �                 �SzH?)�5�	��?       p�C7�R@@�       �                  PV��?�]
���?       ��Ј�7@�       �                 ��%�?$ k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?�       �                    �?��Q#p�?	       ���-3@������������������������       �               H�4H�4@�       �                  c
8?$��C/��?       �~*@�       �                  `�J�?Hy��]0�?       ���y"(@�       �                 ���?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0#@������������������������       �      ��       H�4H�4@������������������������       �      �<       ��#���?�       �                 @  �?�;[��G�?       �O�;�]!@������������������������       �      �<       ���-��@�       �                 �fQ?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 ��C�?8w�;B��?       ՟���	0@������������������������       �        
       �C=�C=,@������������������������       �      ȼ       ��/����?�       �                 �=�t?l���W�?E       �gZSL_@�       �                 P<�\?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 `�0z? $OA�?C       P�v��^@�       �                 ���o?��¡�r�?       �'��!�:@�       �                 ��f?l*�'=P�?        �22@������������������������       �               ��/����?�       �                  s��?�6��b�?       &�|�1@������������������������       �               ��/����?������������������������       �               0#0#0@�       �                 @*��?�;[��G�?       �O�;�]!@������������������������       �               0#0#�?������������������������       �      ��       ��/���@�       �                 P!d�?��Q]K��?6       F�_�W@������������������������       �               ��+��+D@�       �                 �bW�?����?       h�j[��K@�       �                  �E�?��;�� �?       ).���4@�       �                  `���?�'z�3�?       ���da�%@�       �                 p�B�?d����?       �����!@������������������������       �      ��       �C=�C=@������������������������       �      �<       ��/����?������������������������       �      ȼ       ��/����?������������������������       �               ��+��+$@�       �                    �?      �<       S2%S2%A@������������������������       �               #0#06@������������������������       �               H�4H�4(@�t�bh�hhK ��h��R�(KK�KK��h �B�  u�}e@�]�ڕ�`@��-��-e@cCy��d@6��18^@�A�AN@���khc@��F:l$Z@H�4H�48@�}��a@F�JԮDQ@%S2%S27@j1��tVQ@���-��J@��)��)3@�P^CyO@F�JԮDA@��+��+$@\Lg1��6@鰑5@0#0#�?;��,��@��On�(@        ��#���?/����/#@                0����/@                ��/����?                ��/���@        ��#���?0����/@        ��#���?                        0����/@        ��#��@�cp>@        ��#�� @                ��#�� @�cp>@                ��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ��,���1@D�JԮD!@0#0#�?;��,��@��/���@        ��#��@                ��#���?��/���@                0����/@        ��#���?�cp>@        ��#���?                        �cp>@        |�5��(@��/����?0#0#�?|�5��(@��/����?        z�5��@                z�5��@��/����?                ��/����?        z�5��@                                0#0#�?������C@���-��*@vb'vb'"@��#��0@鰑%@H�4H�4@                0#0#@��#��0@鰑%@0#0# @��#��0@���-��@0#0# @��#���?�cp>@0#0#�?��#���?        0#0#�?��#���?                                0#0#�?        �cp>@        �P^Cy/@��/���@0#0#�?        ��/����?        �P^Cy/@�cp>@0#0#�?�P^Cy/@�cp>@        �k(��"@�cp>@        �k(��"@��/����?        �k(��"@                        ��/����?                ��/����?        z�5��@                                0#0#�?        ��/���@                ��/����?                �cp>@        [Lg1��6@�cp>@H�4H�4@[Lg1��6@��/����?0#0# @\Lg1��6@��/����?0#0# @                0#0# @ZLg1��6@��/����?        ��#�� @��/����?        z�5��@                ��#�� @��/����?                ��/����?        ��#�� @                ���>��,@                        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?���>��@0����/3@vb'vb'"@��#��@/����/3@vb'vb'"@��#���?��On�(@        ��#���?0����/@        ��#���?                        0����/@                ��/���@        z�5��@���-��@vb'vb'"@                H�4H�4@z�5��@���-��@H�4H�4@��#���?���-��@        ��#���?��/����?        ��#���?                        ��/����?                0����/@        ��#�� @        H�4H�4@                H�4H�4@��#�� @                z�5��@                ��#���?                ��#�� @                �k(��R@��/���.@0#0#@�P^CyO@��/���@        ��#���?��/����?        ��#���?                        ��/����?        ��>���N@�cp>@        �>��nK@�cp>@        ��#��@@��/����?        �P^Cy?@                ��#�� @��/����?        ��#�� @                        ��/����?        �k(���5@0����/@                ��/����?        �k(���5@�cp>@        �k(��2@��/����?        ���>��,@                ��#��@��/����?        ��#��@                        ��/����?        z�5��@��/����?        ��#�� @                ��#���?��/����?                ��/����?        ��#���?                z�5��@                {�5��(@��/���@0#0#@        0����/@0#0# @        0����/@                        0#0# @|�5��(@�cp>@0#0# @<��,��$@                ��#�� @�cp>@0#0# @��#���?�cp>@0#0# @��#���?�cp>@                ��/����?        ��#���?��/����?        ��#���?                        ��/����?                        0#0# @��#���?                [Lg1��&@����z�A@0#0#�?[Lg1��&@0����/3@0#0#�?��#���?�cp>'@                E�JԮD!@        ��#���?�cp>@        ��#���?                        �cp>@        <��,��$@��/���@0#0#�?                0#0#�?;��,��$@��/���@        ��#���?��/���@                ��/���@        ��#���?                �k(��"@��/���@        ��#��@�cp>@                ��/����?        ��#��@��/����?        z�5��@                ��#���?��/����?                ��/����?        ��#���?                ;��,��@��/����?        ;��,��@                        ��/����?                Nn��O0@                �cp>@                ���-��*@        z�5��(@Nn��O0@vb'vb'B@z�5��(@��|��,@#0#06@<��,��$@��/����?��+��+@                0#0#@;��,��$@��/����?0#0#�?;��,��$@        0#0#�?                0#0#�?<��,��$@                        ��/����?        ��#�� @���-��*@S2%S2%1@��#�� @�cp>@0#0#0@��#���?��/���@                ��/���@        ��#���?                ��#���?��/����?0#0#0@                H�4H�4@��#���?��/����?��+��+$@        ��/����?��+��+$@        ��/����?0#0#@        ��/����?                        0#0#@                H�4H�4@��#���?                        ��/���@0#0#�?        ���-��@                ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?�C=�C=,@                �C=�C=,@        ��/����?        ��#���?��|��,@�;�;[@��#���?��/����?        ��#���?                        ��/����?                ���-��*@�;�;[@        0����/#@S2%S2%1@        ��/����?0#0#0@        ��/����?                ��/����?0#0#0@        ��/����?                        0#0#0@        ��/���@0#0#�?                0#0#�?        ��/���@                ��/���@�q��V@                ��+��+D@        ��/���@|˷|˷I@        ��/���@S2%S2%1@        ��/���@�C=�C=@        ��/����?�C=�C=@                �C=�C=@        ��/����?                ��/����?                        ��+��+$@                S2%S2%A@                #0#06@                H�4H�4(@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJpVhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK煔h��B�2         �                 ���b?Q0�T�?+      G����}@       �                 �H�?s����;�?�       T�{�g?w@       �                 �6��?�lw�K�?�       �5Q�r@       _                 0vb�?�2r��[�?�       a�]�?�n@       ^                  �p�?�CȋS��?f       �H~`"d@       S                 p�v�?�>T����?d       �^x_v@c@       :                  �F�?[f�]e�?V       d ��{�`@                         `��?
UO~��?A       �(qxZ@	       
                 X��>?�`@s'��?       Ei_y,*@������������������������       �               ��#���?������������������������       �               �cp>@                        ��R?�;&����?=       [ɒD��X@                         �^��?Fͻ�&��?       |���g�1@                        �U�?�L����?	       Zk���>)@                         Pmj�?
4=�%�?       �(J��@������������������������       �               ��#�� @������������������������       �               �cp>@                        h��?      �<       ��/���@������������������������       �               ��/����?������������������������       �               �cp>@������������������������       �      �<       ;��,��@                        0��?����?2       ;�nN�RT@������������������������       �               ��/����?       /                 �Y��?�o����?1       ���V��S@                        �<��>��H\i1�?         �?���J@                        �Y�j?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @                        P��?���:z{�?       z��F�H@������������������������       �               ��b:��*@       .                 -��?X����?       ��x��A@        )                 �U����x�<�?       Y&b��qA@!       (                 �Y�b?�����?       �Ä�>c(@"       #                �O�)?`n����?       ~��Y-"@������������������������       �               ��/����?$       %                 hs5�?����?       ��X�)B @������������������������       �               z�5��@&       '                 xi(T?�Z�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@������������������������       �               z�5��@*       -                  ����?�(1k��?       �ꁞ9�6@+       ,                 ���m?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@������������������������       �      ��       �k(��2@������������������������       �      �<       ��/����?0       9                  eX�?�Ƙ���?       ����C:@1       8                 �:W>?�KĈ�?       y�Zc�2@2       3                 𕷋?��?	       ��l}�'*@������������������������       �               ��#��@4       5                 �bS?8�c3���?       �uk��!@������������������������       �               �cp>@6       7                 |$j?^n����?       � ��w<@������������������������       �               ��#��@������������������������       �      �<       ��/����?������������������������       �               �cp>@������������������������       �               ���>��@;       N                 pr��?bꖷh�?       c��=@<       E                 @}L�?Dm�u[U�?       �4���5@=       D                   ��?���mf�?       寠�?b#@>       A                 p�?l?�;[��G�?       �O�;�]!@?       @                 �.�\?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?B       C                    �?      �<       �cp>@������������������������       �               �cp>@������������������������       �               �cp>@������������������������       �               0#0#�?F       I                 �HX?Ƴ�F�M�?       S��ڭQ(@G       H                �r ?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@J       M                 ��?a�ox��?       
c��0 @K       L                 ��j?      �<       �C=�C=@������������������������       �               0#0# @������������������������       �               ��+��+@������������������������       �               ��#���?O       R                 �j%?��r{��?       e�6� @P       Q                 p���?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �               0����/@T       [                 �7z?�FS�5�?       ��9Շ2@U       V                  P���?p���A�?
       0gX\-@������������������������       �               /����/#@W       X                 �Hl�?4=�%�?       �(J��@������������������������       �               �cp>@Y       Z                    �?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?\       ]                 �y��?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      ��       �C=�C=@`       y                 _5?f�6P$g�?2       ��d�QU@a       t                 ��? ���/!�?!       6A���(L@b       s                 ����?(_蹽�?       �Ǣ�9H@c       d                � n�_?��v^�n�?       ��m�G@������������������������       �               ��/����?e       r                 ��n�?P�j���?       �HI�G@f       m                  ���?����X��?       (��֞F@g       j                 ��s?ƃ��̧?       (jW�v%D@h       i                  Ц6�?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@k       l                 NK�X?      �<       �YLg1B@������������������������       �        
       ��,���1@������������������������       �               �k(��2@n       o                 ���? 4=�%�?       �(J��@������������������������       �               ��#���?p       q                 p�L�?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �      �<       ��/����?������������������������       �      �<       ��/����?u       v                 �\��?`�z���?       p���f @������������������������       �               z�5��@w       x                �٬Ӌ?    ��?       "F�b@������������������������       �               H�4H�4@������������������������       �               ��#�� @z       {                  ��j?�c����?       ����<@������������������������       �               ;��,��@|       }                 PTϛ?�4��v�?       �Y-"�7@������������������������       �               0����/#@~                        ��N�?�_�A�?	       肵�e`,@������������������������       �               ;��,��@�       �                 0�2�?� �_rK�?       J�@��"@������������������������       �      ��       ��/���@������������������������       �               ;��,��@�       �                 �!�?)����?'       *��UL@�       �                  �x��?n�hn���?        ��E��F@�       �                  �?�Ș���?       �̨	�>4@�       �                 �{N?����o�?       ]���v<3@������������������������       �        	       �cp>'@�       �                 �yQ?xLU���?       h�ҹ^�@������������������������       �               0#0#�?������������������������       �               ���-��@������������������������       �               0#0#�?�       �                 ��Ɩ?4b
y�	�?       P/㔐k9@�       �                 �m��?ؐV0ߵ�?       %�4�r\3@�       �                  `%+�?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                  �P�?p�i�@M�?
       ���wzb0@�       �                 pU�L?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?�       �                 h��1?      �<       ��On�(@������������������������       �               E�JԮD!@������������������������       �               ��/���@�       �                 ���?ln����?       � ��w<@������������������������       �               ��#��@������������������������       �      �<       ��/����?�       �                  �g<�?�<;�`(�?       ��^�&@������������������������       �               ��#��@�       �                    �?�w��d��?       �0���s@������������������������       �               0#0# @�       �                 �K��?���mf�?       毠�?b@������������������������       �               0#0#�?������������������������       �      �<       ��/���@�       �                 0���?��U�T�?'       .�	[<Q@�       �                 U��?z2���?       Z�n��I@������������������������       �               �cp>@�       �                  �a�?��z��?       �h��G@�       �                 pE��?�Y�)��?       `�e @������������������������       �               z�5��@�       �                    �?lutee�?       Q9��@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                  h��?�n���k�?       �-]ƗC@������������������������       �               ��/����?�       �                    �?(L�0�h�?       l�e�C@�       �                 0vb�?��E�B��?
       dߞKC.@������������������������       �               ��+��+$@�       �                 ��]�?hutee�?       Q9��@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                  �x��?      �<       %S2%S27@������������������������       �               0#0# @������������������������       �               ��-��-5@�       �                 H�`�?��"��b�?
       _���d�2@�       �                    �?�����?       ��X�)B @�       �                 �6AH?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �      �<       ;��,��@�       �                 pm��?������?       +�ǟf%@������������������������       �               ��/���@������������������������       �               H�4H�4@�       �                 �Q�?袰@��?E       �<��Y@�       �                 �מ�?t.R�4�?        ^vE�~F@�       �                 �>�?���d��?
       ��GQ�-@�       �                 ��F�?Hy��]0�?       ���y"@������������������������       �               ��+��+@������������������������       �      ȼ       ��/����?�       �                 �٠r?�� ��?       U?
@�!@������������������������       �               �cp>@�       �                    �?z�G���?       '5L�`�@������������������������       �               0#0# @�       �                 �1��?�@G���?       hu��@������������������������       �               0#0#�?�       �                 �B��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?�       �                 ��Ǽ?��v}�?       ���5>@������������������������       �      ��       #0#06@�       �                 @�	�?w�;B��?       ՟���	 @������������������������       �               ��/����?������������������������       �               �C=�C=@�       �                    �?�����?%       j�j[��K@������������������������       �               0#0#0@�       �                 ��{?�&��գ�?       PHYCz�C@�       �                 `�D�?|�G���?       ��%�|@������������������������       �               ��/����?�       �                 ���?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                  �!�?��M��b�?       8��0��A@�       �                 @W�?      �<       ��-��-5@������������������������       �               0#0# @������������������������       �               ��)��)3@�       �                 ���?H�ih�<�?	       ��
,@������������������������       �               ��/����?�       �                 0���?�n���k�?       3��&�*@������������������������       �               �C=�C=@�       �                 ���?Hy��]0�?       ���y"@�       �                 ��I�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0#@�t�bh�hhK ��h��R�(KK�KK��h �B�  �>��d@鰑Nc@������c@�>��d@����-�a@S2%S2%Q@C����b@����/k_@��8��8:@��tӹa@�H��tXU@��)��)3@�b:���S@Rn��OP@0#0#0@�b:���S@Qn��OP@vb'vb'"@B����R@p��F:lI@vb'vb'"@��,���Q@����z�A@        ��#���?�cp>@        ��#���?                        �cp>@        k1��tVQ@�_��e�=@        ���>��@鰑%@        ��#�� @鰑%@        ��#�� @�cp>@        ��#�� @                        �cp>@                ��/���@                ��/����?                �cp>@        ;��,��@                �P^CyO@0����/3@                ��/����?        �P^CyO@D�JԮD1@        ����JG@���-��@        ��#�� @��/����?                ��/����?        ��#�� @                �GpAF@0����/@        ��b:��*@                �P^Cy?@0����/@        �P^Cy?@��/���@        �k(��"@�cp>@        z�5��@�cp>@                ��/����?        z�5��@��/����?        z�5��@                z�5��@��/����?                ��/����?        z�5��@                z�5��@                �k(���5@��/����?        z�5��@��/����?                ��/����?        z�5��@                �k(��2@                        ��/����?        �P^Cy/@鰑%@        ��#�� @鰑%@        ��#�� @0����/@        ��#��@                ��#��@0����/@                �cp>@        ��#��@��/����?        ��#��@                        ��/����?                �cp>@        ���>��@                ;��,��@��/���.@vb'vb'"@��#��@E�JԮD!@vb'vb'"@        ��/���@0#0# @        ��/���@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@                �cp>@                �cp>@                        0#0#�?��#��@��/����?�C=�C=@z�5��@��/����?                ��/����?        z�5��@                ��#���?        �C=�C=@                �C=�C=@                0#0# @                ��+��+@��#���?                ��#���?���-��@        ��#���?��/����?                ��/����?        ��#���?                        0����/@        ��#��@��|��,@        ��#�� @��On�(@                /����/#@        ��#�� @�cp>@                �cp>@        ��#�� @                ��#���?                ��#���?                ��#�� @��/����?        ��#�� @                        ��/����?                        �C=�C=@�P^CyO@&jW�v%4@H�4H�4@����JG@���-��@H�4H�4@=��,��D@���-��@        >��,��D@�cp>@                ��/����?        =��,��D@0����/@        =��,��D@��/���@        ������C@��/����?        z�5��@��/����?                ��/����?        z�5��@                �YLg1B@                ��,���1@                �k(��2@                ��#�� @�cp>@        ��#���?                ��#���?�cp>@        ��#���?                        �cp>@                ��/����?                ��/����?        ;��,��@        H�4H�4@z�5��@                ��#�� @        H�4H�4@                H�4H�4@��#�� @                �P^Cy/@���-��*@        ;��,��@                ;��,��$@���-��*@                0����/#@        ;��,��$@��/���@        ;��,��@                ;��,��@��/���@                ��/���@        ;��,��@                �k(��"@%jW�v%D@�C=�C=@;��,��@<l��F:B@0#0#@        :l��F:2@0#0# @        :l��F:2@0#0#�?        �cp>'@                ���-��@0#0#�?                0#0#�?        ���-��@                        0#0#�?;��,��@9l��F:2@0#0# @��#���?On��O0@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @��#���?��/���.@        ��#���?�cp>@                �cp>@        ��#���?                        ��On�(@                E�JԮD!@                ��/���@        ��#��@��/����?        ��#��@                        ��/����?        ��#��@��/���@H�4H�4@��#��@                        ��/���@H�4H�4@                0#0# @        ��/���@0#0#�?                0#0#�?        ��/���@        �k(��"@E�JԮD1@��-��-E@z�5��@��/���@������C@        �cp>@        z�5��@0����/@������C@z�5��@��/����?H�4H�4@z�5��@                        ��/����?H�4H�4@        ��/����?                        H�4H�4@        �cp>@wb'vb'B@        ��/����?                ��/����?vb'vb'B@        ��/����?��8��8*@                ��+��+$@        ��/����?H�4H�4@        ��/����?                        H�4H�4@                %S2%S27@                0#0# @                ��-��-5@z�5��@/����/#@H�4H�4@z�5��@��/����?        ��#���?��/����?                ��/����?        ��#���?                ;��,��@                        ��/���@H�4H�4@        ��/���@                        H�4H�4@        �cp>'@#0#0V@        ��/���@�z��z�B@        ���-��@0#0# @        ��/����?��+��+@                ��+��+@        ��/����?                �cp>@H�4H�4@        �cp>@                �cp>@H�4H�4@                0#0# @        �cp>@0#0#�?                0#0#�?        �cp>@                ��/����?                ��/����?                ��/����?�s?�s?=@                #0#06@        ��/����?�C=�C=@        ��/����?                        �C=�C=@        ��/���@�˷|˷I@                0#0#0@        ��/���@fJ�dJ�A@        ��/����?0#0# @        ��/����?                ��/����?0#0# @        ��/����?                        0#0# @        ��/����?B�A�@@                ��-��-5@                0#0# @                ��)��)3@        ��/����?H�4H�4(@        ��/����?                ��/����?H�4H�4(@                �C=�C=@        ��/����?��+��+@        ��/����?0#0#�?                0#0#�?        ��/����?                        0#0#@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK߅�h��B�0         �                 ���b?@
s�I�?9      >_Z���}@       �                 ��??5��[���?�       tL<�Q�v@       �                 �W�?"���?�       ����q@       �                 @���?�2�x�?�       ��x��p@       T                  ���?[��39��?�       �%2.��n@       M                 �^Ҧ?�꟒���?{       �0�[p�f@       F                  .:q?jUw~J��?s       �%�cLee@       A                  #�_?�ֿ�[A�?[       +��Vga@	       :                 �`ğ?0�I���?S       A*��Z�_@
                        �j�%?V����?E       ϻ��)Y@                        ,*����@US�?       �g�l�9@                          �P�?
4=�%�?       �(J��@������������������������       �               ��#�� @������������������������       �               �cp>@                           �?�#�Ѵ�?       �)�B�4@������������������������       �        
       ��b:��*@                        �4U�>h����?       P	K��@������������������������       �               z�5��@                        ��T5?����?       ��X�)B@������������������������       �      ��       z�5��@������������������������       �      �<       ��/����?       )                 �T�|?!���6��?2       5���R@       &                 ��l?N�t���?       �o�go�C@       #                 @F���w"T�?       �W����5@                        0�G?���3�g�?       ص5��2@                        ���2?�L����?	       Yk���>)@                        �U�?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      ��       D�JԮD!@       "                 ��Q�?\n����?       � ��w<@        !                 �bY?      �<       ��#��@������������������������       �               ��#�� @������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?$       %                 (�&R?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ��#�� @'       (                 ��C�?��:V��?	       �GP�1@������������������������       �               ��#��0@������������������������       �      �<       ��/����?*       7                  y��?���쁏�?       x��ձ�A@+       4                 @}L�?�ѭ}��?       |q��:@,       1                 Pa��?h��Y C�?       ?��t��7@-       .                  ���?�Tu��?       ����.@������������������������       �      ��	       ���-��*@/       0                 ��{�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?2       3                 8LSR? ����?       ��X�)B @������������������������       �               ��/����?������������������������       �      �<       z�5��@5       6                    �?~��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @8       9                  ���?��j���?       ���z"@������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?;       <                  ��?87uV��?       m}�'�:@������������������������       �        
       ;��,��4@=       @                  ���?�����?       �O��@>       ?                    �?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      ��       z�5��@B       E                 `�.8?��fm���?       �0��z'@C       D                 ���D? ܜ�x�?       d��إV#@������������������������       �               ��#���?������������������������       �      ��       E�JԮD!@������������������������       �               ��#�� @G       J                 P��^?������?       8nҟ��?@H       I                 0;��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?K       L                  9�>��F¯?       �:.�=@������������������������       �               ��/����?������������������������       �               ���>��<@N       S                 ��jm?^��mf�?       寠�?b#@O       P                 `O~�?|�G���?       ��%�|@������������������������       �               0#0#�?Q       R                  �a�?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?������������������������       �      ��       �cp>@U       �                 @�P�?8lm��R�?)       ��g��P@V       g                  �a�?��A�U1�?$       m�q#N@W       X                 P��r?f����m�?       t�VVk?<@������������������������       �               ���-��@Y       f                 0�� ?�C@0�?       �G��C�5@Z       [                 @b�T?�~�Hs=�?
       ��?Z[0@������������������������       �               ��/����?\       a                 `(��?*DG�?	       �ˠ���.@]       `                 0�e�?p�6L�n�?       �E#��h @^       _                 �j�?bn����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               ;��,��@b       e                ��ߜ?��h��?       S�D'�@c       d                 0���?�|2N��?       �3K}@������������������������       �               z�5��@������������������������       �               0#0# @������������������������       �               ��#�� @������������������������       �               ;��,��@h       q                 0vb�?�骄��?       `(����?@i       p                   ҏ�?��]ۀ��?	       F���O(@j       o                 `��?�@����?       ���a�#@k       l                 J���?�� ��?       rp� k@������������������������       �               ��/����?m       n                 �5W�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       �C=�C=@������������������������       �               ��#�� @r       {                 ���?:.as���?       <�J�2�3@s       z                 �z�?��I@�?       �2d�%@t       u                 �?Pw?$ k�Lj�?       �q��l}#@������������������������       �               ��#���?v       y                 8��?�(���?       y��uk!@w       x                 @GH�?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               0����/@������������������������       �      �<       ��#���?|                        P��?l����?       �����!@}       ~                 0���?�v�;B��?       ՟���	 @������������������������       �               ��/����?������������������������       �               �C=�C=@������������������������       �      ȼ       ��/����?�       �                 ���?���`p��?       �����@������������������������       �               0#0#�?�       �                    �?lutee�?       Q9��@������������������������       �               0#0# @�       �                 �=��?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?�       �                  pm�?���:y�?       7��7@������������������������       �               ��/����?�       �                 �<�?�yo�z�?       A"�-V*6@�       �                    �?���!��?       �@��&@������������������������       �               ��/����?�       �                8�{��?�D�-,�?       �D'ŰO@������������������������       �               ��+��+@������������������������       �               ��#���?������������������������       �               �A�A.@�       �                 �w\�?�\�F�M�?       ��ޚ�&@������������������������       �               ��/����?������������������������       �               ��+��+$@�       �                  �X?;�$���?5       ԥ�~.T@�       �                 ���m?�����?       �O��@�       �                 ���g?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      �<       z�5��@�       �                  �{��?v|�?��?1       h�D[ޥR@�       �                 p"��?\��M��?.       ;�/"cQ@�       �                  ����?p>���Z�?       ]�0�5/8@������������������������       �        	       D�JԮD1@�       �                 p��?��Z�ܙ�?       c����@�       �                    �?�@G���?       hu��@�       �                 (�!�?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��/����?�       �                  �6�?^n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?�       �                 p?U�?Z��T'�?        Fuk���F@�       �                  Z�?�Ϭx���?       �"~���@@�       �                 ����?A�f�?g�?       �� ���=@�       �                 ���?p�r{��?       e�6� @�       �                 ���?      �<       �cp>@������������������������       �               ��/����?������������������������       �               0����/@�       �                 X��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 �n�?��o��^�?       PjO���5@�       �                 ��C?�Yj��}�?       ����=.@�       �                 (���?L� P?)�?       ����x�@������������������������       �               ��#��@������������������������       �               0#0#�?�       �                 �΂�?���/��?       5��o��#@�       �                 tpx?2�c3���?       �uk��!@������������������������       �               z�5��@�       �                 ���?r@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@������������������������       �      ܼ       ��#���?�       �                 �9��?�`@s'��?       Ei_y,*@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               ��#��@�       �                   p��?�>s{Ab�?       `I��n'@������������������������       �               鰑%@������������������������       �               0#0#�?�       �                 ����?     ��<       ��+��+@������������������������       �               0#0# @������������������������       �               H�4H�4@�       �                 ��<{? ����<�?K       PKx���[@������������������������       �               ��#�� @�       �                 p�?ěnd��?J       
�X�>I[@�       �                 ���?�'z�3�?       ���da�5@������������������������       �               #0#0&@�       �                 P�!z?������?       +�ǟf%@������������������������       �               H�4H�4@������������������������       �      ��       ��/���@�       �                 �\��?�<��?=       �4�f�U@�       �                 ����?Xo��?�?       �>���~C@�       �                 ��a�?�BE����?       ~�R��3@�       �                  PV��?X�ih�<�?
       ��
,@������������������������       �               ��/����?������������������������       �        	       H�4H�4(@�       �                 hs5�?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �               0����/@�       �                 P�З?      �<       ��)��)3@������������������������       �               0#0#�?������������������������       �               vb'vb'2@�       �                 ����? 0��?#       �*`.7.H@�       �                 �Z�?���fņ�?       ҋ�'8@������������������������       �               %S2%S27@������������������������       �      �<       ��/����?������������������������       �               H�4H�48@�t�b�$     h�hhK ��h��R�(KK�KK��h �B�  ��P^CYe@Y<�œb@������c@u�}e@o>�c0`@Q��N��O@�5��P>b@j
���S@�+��+�K@�5��P>b@������S@;�;�F@�YLg1b@2����/S@k�6k�69@��>���^@\�v%jWK@0#0#@��>���^@��h
�G@0#0# @���W@�'�xr�F@0#0# @�GpAV@=l��F:B@0#0# @%�}��O@����z�A@0#0# @�k(���5@��/���@        ��#�� @�cp>@        ��#�� @                        �cp>@        ������3@��/����?        ��b:��*@                z�5��@��/����?        z�5��@                z�5��@��/����?        z�5��@                        ��/����?        =��,��D@�]�ڕ�?@0#0# @�#���9@���-��*@        �k(��"@��On�(@        z�5��@��On�(@        ��#�� @鰑%@        ��#�� @��/����?        ��#�� @                        ��/����?                D�JԮD!@        ��#��@��/����?        ��#��@                ��#�� @                ��#�� @                        ��/����?        z�5��@                ��#���?                ��#�� @                ��#��0@��/����?        ��#��0@                        ��/����?        �P^Cy/@;l��F:2@0#0# @���>��@E�JԮD1@0#0# @���>��@On��O0@        ��#���?��|��,@                ���-��*@        ��#���?��/����?        ��#���?                        ��/����?        z�5��@��/����?                ��/����?        z�5��@                        ��/����?0#0# @        ��/����?                        0#0# @��#�� @��/����?        ��#�� @                        ��/����?        �#���9@��/����?        ;��,��4@                ;��,��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        z�5��@                z�5��@D�JԮD!@        ��#���?E�JԮD!@        ��#���?                        E�JԮD!@        ��#�� @                Lp�}>@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ���>��<@��/����?                ��/����?        ���>��<@                        ��/���@0#0# @        ��/����?0#0# @                0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@        [Lg1��6@h
��6@��-��-5@\Lg1��6@%jW�v%4@S2%S2%1@��,���1@E�JԮD!@0#0# @        ���-��@        ��,���1@��/����?0#0# @|�5��(@��/����?0#0# @        ��/����?        z�5��(@��/����?0#0# @���>��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ;��,��@                ;��,��@        0#0# @z�5��@        0#0# @z�5��@                                0#0# @��#�� @                ;��,��@                ;��,��@�cp>'@�A�A.@��#�� @��/����?0#0# @        ��/����?0#0# @        ��/����?0#0#�?        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?                �C=�C=@��#�� @                z�5��@0����/#@�C=�C=@z�5��@��/���@        ��#�� @��/���@        ��#���?                ��#���?��/���@        ��#���?�cp>@        ��#���?                        �cp>@                0����/@        ��#���?                        ��/����?�C=�C=@        ��/����?�C=�C=@        ��/����?                        �C=�C=@        ��/����?                ��/����?0#0#@                0#0#�?        ��/����?H�4H�4@                0#0# @        ��/����?0#0#�?        ��/����?                        0#0#�?��#���?��/����?��+��+4@        ��/����?        ��#���?��/����?��+��+4@��#���?��/����?��+��+@        ��/����?        ��#���?        ��+��+@                ��+��+@��#���?                                �A�A.@        ��/����?��+��+$@        ��/����?                        ��+��+$@\Lg1��6@��On�H@0#0# @;��,��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        z�5��@                ��,���1@{%jW�vH@0#0# @��,���1@z%jW�vH@H�4H�4@��#�� @鰑5@0#0#�?        D�JԮD1@        ��#�� @��/���@0#0#�?        �cp>@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        �P^Cy/@�a#6�;@0#0# @�P^Cy/@D�JԮD1@0#0#�?\Lg1��&@D�JԮD1@0#0#�?��#���?���-��@                �cp>@                ��/����?                0����/@        ��#���?��/����?                ��/����?        ��#���?                <��,��$@鰑%@0#0#�?�k(��"@0����/@0#0#�?��#��@        0#0#�?��#��@                                0#0#�?;��,��@0����/@        ��#��@0����/@        z�5��@                ��#���?0����/@        ��#���?                        0����/@        ��#���?                ��#���?�cp>@        ��#���?                        �cp>@        ��#��@                        鰑%@0#0#�?        鰑%@                        0#0#�?                ��+��+@                0#0# @                H�4H�4@��#�� @��/���.@2��-�rW@��#�� @                        ��/���.@2��-�rW@        ��/���@�C=�C=,@                #0#0&@        ��/���@H�4H�4@                H�4H�4@        ��/���@                ��/���@�6k�6�S@        ���-��@0#0#@@        ���-��@��8��8*@        ��/����?H�4H�4(@        ��/����?                        H�4H�4(@        0����/@0#0#�?                0#0#�?        0����/@                        ��)��)3@                0#0#�?                vb'vb'2@        ��/����?7k�6k�G@        ��/����?%S2%S27@                %S2%S27@        ��/����?                        H�4H�48@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��nhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKㅔh��B�1         h                 �M�?%����F�?,      {�0�n}@       M                 `��?W���$d�?�       ��G�k@       <                 �:W>?��o�?s       h�*`�e@       )                 �U���$l̅X��?V        h�3B`@                        pF�T?$�k0at�?8       �d&͇�U@                         .:q?�(���?       �� �0!:@       
                 �㐢?�#�8b�?       �Ǣ�98@       	                  �ǽ>      �<       �cp>7@������������������������       �               ��/����?������������������������       �               h
��6@������������������������       �      �<       ��#���?                        `焘?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?                        �&d?�'��fr�?(       �w�M@                        ��Yd?jQ��?       �s�=�!@������������������������       �               ��#���?                         �P��?h�r{��?       e�6� @                        �I?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ȼ       �cp>@       (                 �N��?��X3��?!       h���I@       #                 �_?�[��YV�?        ���I@                        `Fe�?��z��?       �T����@@                         �Q�?�ʈD��?       �
��
�5@                        ���?N� P?)�?       ����x�$@������������������������       �               ��#�� @������������������������       �               0#0# @������������������������       �               [Lg1��&@       "                  �Q�? ��<��?       t=�x�(@        !                 �B�q?l@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@������������������������       �               z�5��@$       '                 `��}?�C=+��?       b��T|0@%       &                 x4��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      �<	       ���>��,@������������������������       �      �<       ��/����?*       7                   �P�?��-�8I�?       ��X5��D@+       ,                 `�լ?��{@��?       ��I�@2@������������������������       �               ;��,��@-       6                 ��R�?��?       ��l}�'*@.       /                 LMc?�d�$���?       �T�f$@������������������������       �               ��/����?0       3                  \�&?p�j���?       ���z"@1       2                 ��R?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?4       5                 ����>      �<       z�5��@������������������������       �               ��#���?������������������������       �               ;��,��@������������������������       �      Լ       �cp>@8       9                 �wb9?�q�Ptܳ?       R�� 5�7@������������������������       �               ������3@:       ;                pbѡ�?�����?       ��X�)B@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?=       F                  �Q�?\�$!��?       �] �w0F@>       C                  �0��?�.:�c�?       
�Ol2 :@?       B                 P<�\?��/Ѷ?       ���
$6@@       A                  `���?d�r{��?       e�6� @������������������������       �               ��#���?������������������������       �               ���-��@������������������������       �        	       ��|��,@D       E                ��^�t?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@G       J                    �?��{@��?       ��I�@2@H       I                 0� K?�b8�Y�?       FJͰ(@������������������������       �               ��/����?������������������������       �      �<       [Lg1��&@K       L                 � �?b%@�"�?       ��[�@������������������������       �      ��       ��/���@������������������������       �               ��#�� @N       a                 �i�?\z��L�?       pVu�1F@O       R                 ��?!�M����?       >���(B@P       Q                 �Ղ?X�ih�<�?       ��
@������������������������       �               ��/����?������������������������       �               H�4H�4@S       `                 x�}?����!�?       T��N=@T       ]                 � �?PG�:">�?       �K��G:@U       Z                  �P�?d�r{��?       �)i@7@V       W                    �?vf�T6|�?
       y,*��P+@������������������������       �               D�JԮD!@X       Y                 �wq�?�Z�	7�?       j~���@������������������������       �               z�5��@������������������������       �      �<       ��/����?[       \                ��ח?      �<       0����/#@������������������������       �               E�JԮD!@������������������������       �               ��/����?^       _                 p	t�?ln����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               H�4H�4@b       c                 ���?����?       �a�E�$ @������������������������       �               0#0#@d       e                 p=�?r�T���?       ��e[�&@������������������������       �               ��#�� @f       g                 �F��?x�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?i       �                 �H�?��L���?�       @h��o@j       �                  �6�?B����?X       �c�G�a@k       �                 @�?Q��y��?+       n�$��R@l       }                  �9��?Za�J5��?       ��dA�G@m       x                 8O�?�˳J���?       �a2ِ�8@n       u                 �lO�?23#܅�?	       ���A�0@o       t                 `�?�?ʔfm���?       �0��z'@p       q                 ���?�ۜ�x�?       d��إV#@������������������������       �      �<       �cp>@r       s                  ���?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               ��#�� @v       w                  �я�?      �<       0����/@������������������������       �               �cp>@������������������������       �               ��/����?y       z                 �ꀵ?�̥Q)�?       �9C�<�@������������������������       �               H�4H�4@{       |                  ��3�?
4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @~       �                 ��K�?�n�gn��?       �E��ss7@       �                 ����?��q�R�?       C}Ԥ@������������������������       �               ��#�� @�       �                 ��?|�G���?       ��%�|@������������������������       �               0#0#�?�       �                 Pl?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 �[�Z?�x�<�?       X&b��q1@�       �                  漸?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 `�T�? k� ѽ?	       �����.@�       �                 ���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       ��b:��*@�       �                 �
�k?�� ��?       �^`X:@�       �                  �?إ�je��?       ��BLGh0@������������������������       �      ��       ��|��,@������������������������       �               0#0# @�       �                 <�?*^�yU�?       ��7�1�#@�       �                 �r�w?x�G���?       '5L�`�@������������������������       �               H�4H�4@������������������������       �               �cp>@������������������������       �               0#0#@�       �                 @F���U�?-       �I=��P@�       �                 ���?�w��d��?	       ��EsЖ4@�       �                 ���?<�a
=�?       ��l��@������������������������       �               0#0#�?�       �                 �b'�?      �<       �cp>@������������������������       �               ��/���@������������������������       �               ��/����?�       �                 ��l�?�Qk��?       ��Th!�+@�       �                 ����?�@����?       ���a�#@�       �                 �~��?d*�'=P�?        �2"@�       �                 ��}?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               ��+��+@������������������������       �      ȼ       ��/����?������������������������       �      �<       ��/���@�       �                 �x�?(�����?$       ������G@�       �                 0���?0�Q��?       ���,c�A@�       �                 ���?��(v��?
       �A�s(.@������������������������       �               H�4H�4(@�       �                  �6��?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                  s��?w����?       ��4@�       �                 �x�?fȃ����?       2�i?�{.@�       �                 ����?�djH�E�?	       `�\m�n(@�       �                 p��?�f@���?       hy���"@������������������������       �               0#0# @������������������������       �      ��       ���>��@�       �                  ���?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               H�4H�4@�       �                 p0��?���mf�?       毠�?b@������������������������       �      �<       ��/���@������������������������       �               0#0#�?�       �                 �x��?      �<	       H�4H�4(@������������������������       �               0#0#�?������������������������       �               #0#0&@�       �                 ��o�?�����?E       8%	xp�[@�       �                 �٠�?�&C�:�?6       ]x;�ìU@�       �                 �-�?�.�)���?%       (�ݧ]�O@�       �                  �g<�?�����?       "�D��F@������������������������       �               �cp>@�       �                  @��?���2sW�?       A_8�	D@�       �                 �fQ?��q-��?       j��e|B@�       �                 �q��?�,�#6?�?       ���*4@�       �                 ؼw�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               vb'vb'2@�       �                 ��?�K����?
       B1��0@�       �                 ���`?$�Jg@��?       ��G� �%@������������������������       �               ��/���@�       �                  /Ա?�AP�9��?       i��6��@�       �                 ��?      �<       ��+��+@������������������������       �               0#0#�?������������������������       �               0#0#@������������������������       �      ȼ       ��/����?������������������������       �               H�4H�4@������������������������       �      �<       z�5��@�       �                 xx^�?�C>�?       �1�m�1@������������������������       �               0#0# @�       �                 �S�Y?Ȕfm���?
       ��Z�N/@�       �                 ���R?4=�%�?        �(J��#@�       �                 ��6�?Ĕfm���?       ��Z�N@�       �                   ��?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ȼ       0����/@������������������������       �               ��#�� @������������������������       �               �cp>@�       �                 h~h�?      �<       %S2%S27@������������������������       �               0#0#�?������������������������       �               #0#06@������������������������       �               k�6k�69@�t�bh�hhK ��h��R�(KK�KK��h �BH  �}��a@�xr�'we@��jc@W^CyeZ@�cp>W@��)��)3@ZUUUU�X@E�JԮDQ@��+��+@cCy��T@鰑E@0#0# @�,����G@;l��F:B@0#0# @z�5��@�cp>7@        ��#���?�cp>7@                �cp>7@                ��/����?                h
��6@        ��#���?                ��#�� @                ��#���?                ��#���?                �GpAF@���-��*@0#0# @��#�� @���-��@        ��#���?                ��#���?���-��@        ��#���?��/����?                ��/����?        ��#���?                        �cp>@        ���#8E@���-��@0#0# @���#8E@�cp>@0#0# @��b:��:@0����/@0#0# @������3@        0#0# @��#�� @        0#0# @��#�� @                                0#0# @[Lg1��&@                ���>��@0����/@        ��#���?0����/@        ��#���?                        0����/@        z�5��@                �P^Cy/@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ���>��,@                        ��/����?        �YLg1B@�cp>@        ��b:��*@0����/@        ;��,��@                ��#�� @0����/@        ��#�� @��/����?                ��/����?        ��#�� @��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        z�5��@                ��#���?                ;��,��@                        �cp>@        \Lg1��6@��/����?        ������3@                z�5��@��/����?        z�5��@                        ��/����?        ���>��,@���-��:@H�4H�4@��#���?h
��6@H�4H�4@��#���?鰑5@        ��#���?���-��@        ��#���?                        ���-��@                ��|��,@                ��/����?H�4H�4@        ��/����?                        H�4H�4@��b:��*@0����/@        ZLg1��&@��/����?                ��/����?        [Lg1��&@                ��#�� @��/���@                ��/���@        ��#�� @                ���>��@�cp>7@�C=�C=,@;��,��@h
��6@vb'vb'"@        ��/����?H�4H�4@        ��/����?                        H�4H�4@;��,��@鰑5@H�4H�4@;��,��@鰑5@        z�5��@%jW�v%4@        z�5��@鰑%@                D�JԮD!@        z�5��@��/����?        z�5��@                        ��/����?                0����/#@                E�JԮD!@                ��/����?        ��#�� @��/����?                ��/����?        ��#�� @                                H�4H�4@��#�� @��/����?��+��+@                0#0#@��#�� @��/����?0#0#�?��#�� @                        ��/����?0#0#�?                0#0#�?        ��/����?        d:��,&C@i
���S@R��N�a@�P^Cy?@�a#6�K@�+��+�K@\Lg1��6@�+Q��B@�C=�C=,@[Lg1��6@%jW�v%4@��+��+@;��,��@On��O0@H�4H�4@z�5��@���-��*@        z�5��@E�JԮD!@        ��#���?D�JԮD!@                �cp>@        ��#���?�cp>@        ��#���?                        �cp>@        ��#�� @                        0����/@                �cp>@                ��/����?        ��#�� @�cp>@H�4H�4@                H�4H�4@��#�� @�cp>@                �cp>@        ��#�� @                ��,���1@��/���@0#0# @��#�� @��/����?0#0# @��#�� @                        ��/����?0#0# @                0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?        �P^Cy/@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ���>��,@��/����?        ��#���?��/����?                ��/����?        ��#���?                ��b:��*@                        D�JԮD1@vb'vb'"@        ��|��,@0#0# @        ��|��,@                        0#0# @        �cp>@�C=�C=@        �cp>@H�4H�4@                H�4H�4@        �cp>@                        0#0#@��#�� @:l��F:2@�ڬ�ڬD@        �cp>'@vb'vb'"@        �cp>@0#0#�?                0#0#�?        �cp>@                ��/���@                ��/����?                �cp>@0#0# @        ��/����?0#0# @        ��/����?0#0# @        ��/����?H�4H�4@        ��/����?                        H�4H�4@                ��+��+@        ��/����?                ��/���@        ��#�� @���-��@0#0#@@��#�� @���-��@��+��+4@        ��/����?�C=�C=,@                H�4H�4(@        ��/����?0#0# @        ��/����?                        0#0# @��#�� @�cp>@H�4H�4@��#�� @��/����?��+��+@��#�� @��/����?0#0# @���>��@        0#0# @                0#0# @���>��@                ��#���?��/����?        ��#���?                        ��/����?                        H�4H�4@        ��/���@0#0#�?        ��/���@                        0#0#�?                H�4H�4(@                0#0#�?                #0#0&@���>��@�e�_��7@��+��+T@���>��@�e�_��7@�+��+�K@���>��@�e�_��7@0#0#@@z�5��@��On�(@�A�A>@        �cp>@        z�5��@���-��@�A�A>@        ���-��@�A�A>@        ��/����?��)��)3@        ��/����?0#0#�?                0#0#�?        ��/����?                        vb'vb'2@        �cp>@#0#0&@        �cp>@��+��+@        ��/���@                ��/����?��+��+@                ��+��+@                0#0#�?                0#0#@        ��/����?                        H�4H�4@z�5��@                ��#��@�cp>'@0#0# @                0#0# @��#��@�cp>'@        ��#��@�cp>@        ��#�� @�cp>@        ��#�� @��/����?                ��/����?        ��#�� @                        0����/@        ��#�� @                        �cp>@                        %S2%S27@                0#0#�?                #0#06@                k�6k�69@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJXk�hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKɅ�h��B�+         �                 �6Sz?GP5�R�?#      bъG7y}@       �                 p���?�t��_�?�       ʱ V�x@       v                 �"��?��Q.;�?�       w� ��Su@       a                 0�{?qv
+���?�       ��踱�o@       H                 P�f�?�����?r       m2Elg@       3                  �v�?f�� H��?X       \<�œb@       &                 `%�7?u��	��?G       ��N0g�]@                         �3��?�g�?� �?2       C~aƍU@	       
                 `f��>΃�\��?       �D+զm7@������������������������       �               ��/����?                         `s�?`����?       �Fx�v�5@                         Џ~�?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?                        p�־?�hK)�?       �h��K�2@������������������������       �               z�5��(@                        ��p?�����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?       %                 ��q?��V���?"       �fX�dO@                         �U���ζ�Ӣ�?       D����J@                        �2*�?�&��$C�?       ���+p8@                        ���?�3+�Pr�?       Z-"�=L4@                        `f��>��|��?       ���ĺw@������������������������       �               0����/@������������������������       �               ��#�� @                        .25Q?      �<       ���-��*@������������������������       �               ��On�(@������������������������       �               ��/����?                        ��cr?      �<       ��#��@������������������������       �               ��#�� @������������������������       �               ��#�� @!       $                 x��?�]���?       �j0�W�<@"       #                   E(�?jP�D�?       �A��P?$@������������������������       �               �cp>@������������������������       �               ���>��@������������������������       �        
       �k(��2@������������������������       �               /����/#@'       2                 Pc	�?3#܅�?       ���A�@@(       1                  0p��?d�r{��?       e�6� ?@)       0                    �?�u�N��?       ������=@*       +                  �~��?�`@s'��?       �[�_4@������������������������       �      ��	       ��On�(@,       -                 ��i?Fǵ3���?       �q�ͨ�@������������������������       �               ��#�� @.       /                 ��[?r@ȱ��?       om���S@������������������������       �               0����/@������������������������       �               ��#���?������������������������       �               0����/#@������������������������       �      �<       ��#���?������������������������       �      �<       ��#�� @4       G                 �Q�?�@US�?       �g�l�9@5       D                    �?��6L�n�?       ��4}i�8@6       A                 �@�?�q���?       ��|�^1@7       >                 �E�+? M�����?	       p����.@8       =                 �-�?h�s�	�?       f���*@9       <                  Џ~�?����?       ��X�)B@:       ;                 ��aӾ���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �               �k(��"@?       @                 �_��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?B       C                  p���?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?E       F                 h��?      �<       ���>��@������������������������       �               ��#���?������������������������       �               z�5��@������������������������       �      �<       ��/����?I       ^                  ��?�\�,�?       <�/ZBE@J       Q                 ��
q?����?       �U0C@K       L                  L��?�AP�9��?       i��6��+@������������������������       �               ��+��+@M       N                    �?�Ϟi�?       
��ؠ�!@������������������������       �               �cp>@O       P                  �0��?Fy��]0�?       ���y"@������������������������       �               ��+��+@������������������������       �      ȼ       ��/����?R       [                 ��^�?�[�*��?       Q��s8@S       X                 �~�?&�g���?       ���u3@T       W                  `���?�@����?       ���a�@U       V                 (o��?z��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               0#0# @Y       Z                 ��li?��&���?
       ��G2��,@������������������������       �               ��#���?������������������������       �        	       ���-��*@\       ]                 �u�y?�@����?       ���a�@������������������������       �               ��/����?������������������������       �               0#0#@_       `                  P���?      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@b       o                  �g<�?���;z�?(       ÀG91�P@c       l                 �C�Z?�B	���?       �$r.X{?@d       k                  ys8?�Z�!���?       ��e`��<@e       f                    �?��?       ��l}�'*@������������������������       �               ��/���@g       j                 �,�?X�j���?       ���z"@h       i                 X�)�?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@������������������������       �               ;��,��@������������������������       �      ��       �P^Cy/@m       n                    �?     ��<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?p       u                 P�?���=l>�?       7�U[��A@q       r                 ԰�C?�Ͳ�S{�?       pս��i3@������������������������       �      �<	       �P^Cy/@s       t                 ,	�?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �               ��#��0@w       |                   ��?������?7       F���˘U@x       {                 ��6�?�^�#΀�?       O�{��A5@y       z                 �ڡ3?      �<
       /����/3@������������������������       �               0����/@������������������������       �               ��|��,@������������������������       �      ܼ       ��#�� @}       �                 �U�<?�̣��B�?,       5�� VHP@~       �                 p-�?ޗ,�!�?       -%�I4�@@       �                 �Q��?�<�Aw��?       8&�+o|(@������������������������       �               ���>��@�       �                ��G��?��b�}�?       ���\�@�       �                  4�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               ��#�� @�       �                 �~��?�Ñp��?       <7��0�5@�       �                    �?�v�;B��?       ՟���	 @������������������������       �               0#0# @�       �                 `Fe�?Hy��]0�?       ���y"@������������������������       �               ��/����?������������������������       �               ��+��+@�       �                 @��?�T�"��?
       ��`2�Z+@�       �                  P�"�?�;[��G�?       �O�;�]!@������������������������       �               ��/���@�       �                 �:�{?���mf�?       毠�?b@������������������������       �               0#0#�?������������������������       �      �<       ��/���@�       �                 �.!�?�@����?       ���a�@������������������������       �               ��/����?������������������������       �               0#0#@�       �                 `�?D��ce�?       z����0?@�       �                 ��`�?L+�P���?       �%�8�3@�       �                 (ww�?���mf�?       寠�?b#@�       �                 @���?�;[��G�?       �O�;�]!@������������������������       �               0#0#�?������������������������       �      �<       ��/���@������������������������       �               0#0#�?�       �                 x9I�?*^�yU�?       ��7�1�#@�       �                 ضm�?~�G���?       '5L�`�@������������������������       �               ��/����?�       �                 �ş�?����|e�?       �z �B�@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?������������������������       �               0#0#@�       �                 `��?�>s{Ab�?       `I��n'@������������������������       �               0#0#�?������������������������       �               鰑%@�       �                 @8�?&d����?       �b��R�I@�       �                 �;�?�it�R��?       ���O@@�       �                 ��?Ğ��n��?       ����5@�       �                 (�A�?ȏBC��?       �WDl��0@������������������������       �               ��#���?�       �                 `�C?���`�?       ��
�Me/@�       �                 �b'�?�y��d��?       �=�0�@������������������������       �               H�4H�4@�       �                pn�ǣ?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @�       �                 ���?�;[��G�?       �O�;�]!@������������������������       �               0#0#�?������������������������       �               ��/���@�       �                 p�!�?      �<       0����/@������������������������       �               ��/����?������������������������       �               ��/���@������������������������       �               #0#0&@�       �                  R��?xL�0�h�?	       l�e�3@�       �                 �D��d*�'=P�?        �2"@�       �                  �~��?����|e�?       �z �B�@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?������������������������       �               ��+��+@�       �                 p ��?      �<       ��+��+$@������������������������       �               0#0# @������������������������       �               0#0# @�       �                  9ר?�w|ۯ��?5       b~����S@�       �                 h��?H�)�n�?       �b�}{.;@������������������������       �               ��)��)3@�       �                  N��?w�;B��?       ՟���	 @������������������������       �               �C=�C=@������������������������       �      ȼ       ��/����?�       �                 @��?      �<"       |˷|˷I@������������������������       �               H�4H�4@������������������������       �        !       F�4H�4H@�t�bh�hhK ��h��R�(KK�KK��h �B�  y�YLGc@�����d@��)��)c@y�YLGc@��-��bd@�i��R@C����b@��z��wb@��-��-E@}�5�wa@�e�_��W@��)��)3@bCy��T@�H��tXU@vb'vb'2@������S@���|�P@        u�}wL@1����-O@        �}�\I@����z�A@        �k(��2@0����/@                ��/����?        �k(��2@�cp>@        ��#���?��/����?        ��#���?                        ��/����?        ��,���1@��/����?        z�5��(@                ;��,��@��/����?        ;��,��@                        ��/����?        ���b:@@��/���>@        ���b:@@鰑5@        z�5��@:l��F:2@        ��#�� @:l��F:2@        ��#�� @0����/@                0����/@        ��#�� @                        ���-��*@                ��On�(@                ��/����?        ��#��@                ��#�� @                ��#�� @                �#���9@�cp>@        ���>��@�cp>@                �cp>@        ���>��@                �k(��2@                        /����/#@        z�5��@���-��:@        ��#��@���-��:@        z�5��@���-��:@        z�5��@E�JԮD1@                ��On�(@        z�5��@0����/@        ��#�� @                ��#���?0����/@                0����/@        ��#���?                        0����/#@        ��#���?                ��#�� @                �k(���5@��/���@        �k(���5@�cp>@        ���>��,@�cp>@        ��b:��*@��/����?        z�5��(@��/����?        z�5��@��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#�� @                �k(��"@                ��#���?��/����?        ��#���?                        ��/����?        ��#���?��/����?        ��#���?                        ��/����?        ���>��@                ��#���?                z�5��@                        ��/����?        ;��,��@0����/3@vb'vb'2@��#���?0����/3@vb'vb'2@        ��/���@��+��+$@                ��+��+@        ��/���@��+��+@        �cp>@                ��/����?��+��+@                ��+��+@        ��/����?        ��#���?��/���.@0#0# @��#���?��|��,@0#0#@        ��/����?0#0#@        ��/����?0#0# @                0#0# @        ��/����?                        0#0# @��#���?���-��*@        ��#���?                        ���-��*@                ��/����?0#0#@        ��/����?                        0#0#@��#��@                ��#���?                z�5��@                .�����K@鰑%@0#0#�?�,����7@��/���@        �,����7@0����/@        ��#�� @0����/@                ��/���@        ��#�� @��/����?        z�5��@��/����?                ��/����?        z�5��@                ;��,��@                �P^Cy/@                        �cp>@                ��/����?                ��/����?        ���b:@@�cp>@0#0#�?�P^Cy/@�cp>@0#0#�?�P^Cy/@                        �cp>@0#0#�?        �cp>@                        0#0#�?��#��0@                [Lg1��&@�cp>�I@%S2%S27@��#�� @/����/3@                /����/3@                0����/@                ��|��,@        ��#�� @                �k(��"@Pn��O@@%S2%S27@�k(��"@�cp>'@��8��8*@�k(��"@��/����?0#0#�?���>��@                ��#�� @��/����?0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?        ��#�� @                        /����/#@H�4H�4(@        ��/����?�C=�C=@                0#0# @        ��/����?��+��+@        ��/����?                        ��+��+@        E�JԮD!@��+��+@        ��/���@0#0#�?        ��/���@                ��/���@0#0#�?                0#0#�?        ��/���@                ��/����?0#0#@        ��/����?                        0#0#@        鰑5@��+��+$@        鰑%@vb'vb'"@        ��/���@0#0# @        ��/���@0#0#�?                0#0#�?        ��/���@                        0#0#�?        �cp>@�C=�C=@        �cp>@H�4H�4@        ��/����?                ��/����?H�4H�4@                H�4H�4@        ��/����?                        0#0#@        鰑%@0#0#�?                0#0#�?        鰑%@        z�5��@��/���.@B�A�@@z�5��@��|��,@�A�A.@z�5��@��|��,@0#0#@z�5��@/����/#@0#0#@��#���?                ��#�� @0����/#@0#0#@��#�� @��/����?H�4H�4@                H�4H�4@��#�� @��/����?                ��/����?        ��#�� @                        ��/���@0#0#�?                0#0#�?        ��/���@                0����/@                ��/����?                ��/���@                        #0#0&@        ��/����?vb'vb'2@        ��/����?0#0# @        ��/����?H�4H�4@                H�4H�4@        ��/����?                        ��+��+@                ��+��+$@                0#0# @                0#0# @        ��/����?��jS@        ��/����?��8��8:@                ��)��)3@        ��/����?�C=�C=@                �C=�C=@        ��/����?                        |˷|˷I@                H�4H�4@                F�4H�4H@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ0��JhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK酔h��B�2         z                  ��d�?��w�T�?'      a�!F�}@       [                 ��H?ԕ��?�       ��)	�l@       N                 pm��?�*���|�?a       ��]d@                          �G�?�}+ǎ��?R       i~u_R�`@                        P]ڒ?b-����?       �T|qt�>@                        ��?��I@�?       �2d�5@                         �[6?� �_rK�?       J�@��"@                           �?<9�)\e�?       _���b @	       
                 ��k?�����?       �O��@������������������������       �               ��/����?������������������������       �      �<       ;��,��@������������������������       �      �<       ��/����?������������������������       �      м       ��/����?                        �M}C?D��c`�?       %��t5)@������������������������       �               �cp>'@������������������������       �      ܼ       ��#���?                         �G?�?L���'0�?       �C�� T"@                          S�?      �<       ;��,��@������������������������       �               ��#���?������������������������       �               ��#��@                        �)�(?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?       3                  �P��?LXO�#�??       �狢G Z@       2                  P��?b��
�?       ���TH@                        P�1?� y�m�?       {��<�G@                           �?�)z� ��?       �\�@                       �(�!?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �      �<       ��/����?        '                 ��T�?6�(��?       ��� �D@!       "                 p`�? ���OT�?       p�>%,�9@������������������������       �      ȼ       ZLg1��6@#       &                    �?dn����?       � ��w<@$       %                 �j%?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#���?(       -                 p�F�?��Fl�R�?
       ��޷/�,@)       ,                   .p�?=�N9���?       ��{j�@*       +                 �ѱ?f,���O�?       ���/>@������������������������       �               ��#���?������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?.       /                 �&p?h�j���?       ���z"@������������������������       �               ��/����?0       1                 ��?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ���>��@������������������������       �     ��<       0#0#�?4       K                 ��x�?�G�&�?"       Է{G:5L@5       F                 @��?�c�ǰ(�?       �^�mƦH@6       ?                 ���?4�^��?       B<��*�B@7       >                 @�>?�q���?       ��|�^1@8       =                 D�C'?�)z� ��?       ��\�@9       :                   �P�?�d�$���?       �T�f@������������������������       �               z�5��@;       <                  L��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      �<       ��/����?������������������������       �               <��,��$@@       E                 `�
E?��|��?       ³�̙4@A       B                 �Y�b?�FS�5�?       ��9Շ2@������������������������       �        	       �cp>'@C       D                 ���?�)z� ��?       �\�@������������������������       �               ��#��@������������������������       �               �cp>@������������������������       �      �<       ��#�� @G       H                 8���?2��/��?       ��t�o�&@������������������������       �               ��#�� @I       J                 p|��?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?L       M                 8���?��3Fi�?       :�"Ξs@������������������������       �               ��+��+@������������������������       �               ��#�� @O       V                 0y��?�zH3�?       +��Z�9@P       U                 `۶�?j��#n�?	       u���/@Q       R                 p;ݩ?8��~d��?       7E���*@������������������������       �               �cp>'@S       T                  �/�?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��#�� @W       Z                    �?Ƣ��'�?       �^��$@X       Y                 �[��?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               �C=�C=@\       ]                 0��?�u�O2�?,       L��V)Q@������������������������       �               E�JԮD!@^       q                  �g<�?:@8)�q�?'       Ha� �N@_       b                 `.�?hV�\Ga�?       q�6tE@`       a                 �i?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@c       d                  ^ߵ?�Zz.��?       �`K�kC@������������������������       �               0#0# @e       p                 ��@p?�F&�u{�?       �0(�iB@f       k                 ��{�?x��OU�?       qp���?@g       h                 Ё��?���mf�?       毠�?b@������������������������       �               �cp>@i       j                  K�V?~�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?l       m                 p��? �m���?       vD���:@������������������������       �               &jW�v%4@n       o                 `TF�?�`@s'��?       Ei_y,*@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               ��+��+@r       u                 ���?����?       ~�5�1@s       t                 ���?L� P?)�?       ����x�@������������������������       �               ��#��@������������������������       �               0#0#�?v       y                 ��C�?����|e�?       8\@��'@w       x                 �+�[?��H�&p�?       L^�3��%@������������������������       �               ��/����?������������������������       �               vb'vb'"@������������������������       �      м       ��/����?{       �                 0��?׶6�C�?�       9�/�Tn@|       �                 �je?*p{��?O       ��Q�Ku_@}       �                 ��(�?8���0�?E       d7I+�l[@~       �                  ���?P�|9��?4       ��Dp��S@       �                  ���+��?       �|��C@�       �                  ����?`n����?       � ��w<(@�       �                    �?� �_rK�?       J�@��"@�       �                 �;�?�d�$���?       �T�f@������������������������       �               z�5��@�       �                 `]j�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 �c�?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �      �<       z�5��@�       �                  �Q�?.�r?�?       �M�)#�;@�       �                  l@?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      �<       �#���9@�       �                  @���?`��ڄy�?       �P�cG�C@�       �                 p۶�?t�a����?       ��� �CB@�       �                 `���?x�\~�s�?       ����y<@�       �                 ��x�?u!\��?       ��\��5@�       �                 p�i?��_�u��?       ��X̰3@������������������������       �               �cp>@�       �                 �_��?�&�+�?       q��wy�+@�       �                 ��ۜ?B�pB}��?       ����1$@�       �                  ���?d����?       Q	K��@�       �                 �-�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               ��#��@�       �                 ����?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �      ��       ��/���@�       �                 �Xx�?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?������������������������       �      ��       ���-��@�       �                 Xi?69�)\e�?       _���b @�       �                 p}<l?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               ��#��@������������������������       �               z�5��@�       �                 �j�?�g}��?       i��>>@�       �                 �HX?��jts^�?
       ��4`,/2@�       �                ��r?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                  ����?a�ox��?       
c��00@������������������������       �               ��#�� @�       �                 ���z?      �<       �C=�C=,@������������������������       �               0#0#@������������������������       �               ��+��+$@�       �                 �j%?B��NV=�?       �W�%�'@�       �                ����?�J���?       a���@������������������������       �               H�4H�4@������������������������       �               z�5��@�       �                  �0��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/���@�       �                    �?      �<
       0#0#0@������������������������       �               H�4H�4@������������������������       �               ��8��8*@�       �                 `}�?�K1+�I�?K       �\}�3]@�       �                 pJ�q?��E$	�?5       �{%i��T@�       �                 ����?�-"�)��?       ���6<B@�       �                 ��{�?:jk�5�?       �R�3A@������������������������       �               H�4H�4@�       �                  0���?���G���?       a]���X<@�       �                 ��?^��Yy��?       lo�D9@�       �                 �H��?|�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 @���?@�+���?       �aJ9U5@�       �                    �?f%@�"�?       �6�E�!@�       �                 �1�?      �<       0����/@������������������������       �               ��/����?������������������������       �               ��/���@�       �                 3��?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@������������������������       �      �<	       ��On�(@�       �                 J;h�?^����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?������������������������       �      �<       ��#�� @�       �                 (F�? xUA�u�?       �W����G@�       �                 �	��?�w��d��?       �0���s@������������������������       �      �<       H�4H�4@������������������������       �               ��/���@�       �                 ��M�?`,�#6?�?       ���*D@�       �                 �Qz�?Hy��]0�?       ���y"@������������������������       �               0#0#@�       �                 Hн�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                    �?�5���?       ��P9�A@������������������������       �      ȼ
       ��)��)3@�       �                 hp�?��(v��?	       �A�s(.@������������������������       �               ��8��8*@�       �                 �>��?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 ����? �;{���?       ���'Ν@@������������������������       �               ��/����?������������������������       �               0#0#@@�t�bh�hhK ��h��R�(KK�KK��h �B�  �>��d@������c@�؉��Ic@�,����W@�œ[<9X@�z��z�B@�k(���U@\�v%jWK@��)��)3@bCy��T@(jW�v%D@#0#0&@��b:��*@E�JԮD1@        z�5��@��/���.@        ;��,��@��/���@        ;��,��@�cp>@        ;��,��@��/����?                ��/����?        ;��,��@                        ��/����?                ��/����?        ��#���?�cp>'@                �cp>'@        ��#���?                ���>��@��/����?        ;��,��@                ��#���?                ��#��@                ��#�� @��/����?        ��#�� @                        ��/����?        ��,���Q@�cp>7@#0#0&@d:��,&C@�cp>@0#0#@d:��,&C@�cp>@H�4H�4@��#��@�cp>@        ��#��@��/����?        ��#��@                        ��/����?                ��/����?        Ey�5A@�cp>@H�4H�4@|�5��8@��/����?        ZLg1��6@                ��#�� @��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#���?                �k(��"@��/����?H�4H�4@��#���?��/����?H�4H�4@��#���?        H�4H�4@��#���?                                H�4H�4@        ��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ��#���?                ���>��@                                0#0#�?���b:@@E�JԮD1@�C=�C=@Jp�}>@E�JԮD1@0#0# @<��,��4@E�JԮD1@        ���>��,@�cp>@        ��#��@�cp>@        ��#��@��/����?        z�5��@                ��#���?��/����?        ��#���?                        ��/����?                ��/����?        <��,��$@                z�5��@��|��,@        ��#��@��|��,@                �cp>'@        ��#��@�cp>@        ��#��@                        �cp>@        ��#�� @                �k(��"@        0#0# @��#�� @                ��#���?        0#0# @                0#0# @��#���?                ��#�� @        ��+��+@                ��+��+@��#�� @                z�5��@��|��,@0#0# @��#�� @��On�(@0#0#�?        ��On�(@0#0#�?        �cp>'@                ��/����?0#0#�?        ��/����?                        0#0#�?��#�� @                ��#���?��/����?�C=�C=@��#���?��/����?        ��#���?                        ��/����?                        �C=�C=@��#�� @鰑E@vb'vb'2@        E�JԮD!@        ��#�� @�-����@@vb'vb'2@��#��@��/���>@0#0# @z�5��@��/����?                ��/����?        z�5��@                ��#���?�_��e�=@0#0# @                0#0# @��#���?�_��e�=@H�4H�4@��#���?�_��e�=@0#0#�?        ��/���@0#0#�?        �cp>@                ��/����?0#0#�?                0#0#�?        ��/����?        ��#���?�cp>�9@                &jW�v%4@        ��#���?�cp>@        ��#���?                        �cp>@                        ��+��+@��#��@�cp>@��+��+$@��#��@        0#0#�?��#��@                                0#0#�?        �cp>@vb'vb'"@        ��/����?vb'vb'"@        ��/����?                        vb'vb'"@        ��/����?        �P^CyMP@<��18N@ t?�s?]@���>��L@�-����@@S2%S2%A@���>��L@�-����@@vb'vb'2@�#���I@���-��:@0#0#�?��,���A@0����/@        ��#�� @��/���@        ;��,��@��/���@        ��#��@��/����?        z�5��@                ��#���?��/����?                ��/����?        ��#���?                ��#���?�cp>@                �cp>@        ��#���?                z�5��@                ��b:��:@��/����?        ��#���?��/����?                ��/����?        ��#���?                �#���9@                ��#��0@h
��6@0#0#�?��b:��*@h
��6@0#0#�?��#�� @/����/3@0#0#�?��#�� @��On�(@0#0#�?z�5��@��On�(@0#0#�?        �cp>@        z�5��@���-��@0#0#�?z�5��@�cp>@0#0#�?z�5��@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ��#��@                        ��/����?0#0#�?                0#0#�?        ��/����?                ��/���@        ��#�� @                ��#���?                ��#���?                        ���-��@        ;��,��@�cp>@        ��#���?�cp>@        ��#���?                        �cp>@        ��#��@                z�5��@                z�5��@���-��@S2%S2%1@z�5��@��/����?�C=�C=,@��#���?��/����?                ��/����?        ��#���?                ��#�� @        �C=�C=,@��#�� @                                �C=�C=,@                0#0#@                ��+��+$@z�5��@�cp>@H�4H�4@z�5��@        H�4H�4@                H�4H�4@z�5��@                        �cp>@                ��/����?                ��/���@                        0#0#0@                H�4H�4@                ��8��8*@���>��@���-��:@�ڬ�ڬT@���>��@�cp>�9@n�6k�6I@���>��@%jW�v%4@vb'vb'"@;��,��@$jW�v%4@vb'vb'"@                H�4H�4@;��,��@&jW�v%4@H�4H�4@z�5��@&jW�v%4@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @z�5��@:l��F:2@        z�5��@�cp>@                0����/@                ��/����?                ��/���@        z�5��@��/����?                ��/����?        z�5��@                        ��On�(@        ��#�� @        0#0#�?��#�� @                                0#0#�?��#�� @                        �cp>@�ڬ�ڬD@        ��/���@H�4H�4@                H�4H�4@        ��/���@                ��/����?��)��)C@        ��/����?��+��+@                0#0#@        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?B�A�@@                ��)��)3@        ��/����?�C=�C=,@                ��8��8*@        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?0#0#@@        ��/����?                        0#0#@@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJڡWhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK텔h��B�3         �                 ��\�?���J�2�?.      ���h}@       Y                 0-3�?Y�UHu�?�       ߭���q@       J                  .:q?B5�m���?       Po��o]i@                         _z_?on�I��?h       �7bXd@                        �@�F?( k�Lj�?       g*�}#<=@                        �I?@9�)\e�?       `���b @                        X�Oq?4=�%�?       �(J��@                        �y���\n����?       � ��w<@	       
                 d��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#���?������������������������       �               ��/����?������������������������       �               z�5��@                        Va�?@H�,.̷?       �J�$r.5@������������������������       �               'jW�v%4@������������������������       �      �<       ��#���?       ;                  p�:?f��<���?S       N���~�`@       ,                 �vs?2�#ShS�?;       ��I���W@       %                 �U���J&Μ�!�?(       D3�\rN@                        �SO?l�Y�`��?       �����8@                          \��?��Z�	7�?	       ���`�$.@                        �5~S?@ǵ3���?       �q�ͨ�@������������������������       �               0����/@������������������������       �               z�5��@                         h��?P����?       P	K��@                           �?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               ��#��@                         �c-?* k�Lj�?       �q��l}#@������������������������       �               ��#���?!       "                  e_?�(���?       y��uk!@������������������������       �               �cp>@#       $                 p��v?b%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?&       '                 (�+0?`��E2ȹ?       ;�f��	B@������������������������       �      �<       �k(���5@(       )                 �B�U?\����?       P	K��,@������������������������       �               \Lg1��&@*       +                 @F�b%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?-       2                 �{��?v/�B���?       1`��:A@.       1                 ���?p�i�@M�?       ���wzb0@/       0                  ���?h�r{��?       e�6� @������������������������       �               ���-��@������������������������       �               ��#���?������������������������       �      ��       E�JԮD!@3       :                 �-�?��`$��?       xn��*2@4       7                  �d�?���_�?       ���e��#@5       6                  ��?�;�a
=�?       ��l��@������������������������       �               �cp>@������������������������       �               0#0#�?8       9                 �j%?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               ��#�� @<       ?                 �&oh?��_�u��?       ��X̰C@=       >                   ���?\����?       P	K��@������������������������       �               ��/����?������������������������       �               z�5��@@       C                  �Ԧ�?��0���?       Є��@@A       B                  `��?��٤ݸ?       ��<5�84@������������������������       �               ��#���?������������������������       �               /����/3@D       I                 x��y?�\U�?       �{����'@E       F                 `f�?���/��?       6��o��#@������������������������       �               ��/����?G       H                 p#��?@9�)\e�?       _���b @������������������������       �               �cp>@������������������������       �               ;��,��@������������������������       �               0#0# @K       L                   �P�?���4��?       ��v�yC@������������������������       �               z�5��8@M       R                  �E�?)�ť��?       [`Il�7,@N       O                &�rq?����]L�?       N66�ͯ@������������������������       �               ��#���?P       Q                   ��?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@S       V                 `�s�?&A����?       4E���_"@T       U                 tS��?,Lj����?       ���T�@������������������������       �               z�5��@������������������������       �               0#0#�?W       X                 h��?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?Z       �                 0�3�?����g��?0       ���'��Q@[       �                 �*/�?s�H�+�?%       !�AZ6�L@\       ]                 @���>b�1l���?        |�+�~H@������������������������       �               ��#���?^       }                 p�~�?���Y��?       2A#.�G@_       p                 ho��?B���ޙ�?       ��~j�B@`       a                 p���?��,����?       V��L7@������������������������       �               0#0# @b       m                 ��Ĳ?�}>D�P�?       �狢G5@c       j                 `Fe�?�5JH���?       �MOI3@d       i                 0�M�?�� ��?       qp� k@e       h                 (�i<?x��`p��?       �����@f       g                 ���?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               0#0#�?������������������������       �               �cp>@k       l                 `U�?      �<       ���-��*@������������������������       �               D�JԮD!@������������������������       �               0����/@n       o                  �~��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?q       r                 ���{?TC6&x�?
       �V�5,@������������������������       �               H�4H�4@s       z                 �@3�?L
wf�x�?       0����(&@t       u                 �6O�?r�G���?       '5L�`�@������������������������       �               ��/����?v       y                 `��?����|e�?       �z �B�@w       x                 @��?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0# @{       |                 @�F�?      �<       ;��,��@������������������������       �               ��#���?������������������������       �               ��#��@~                           �?      �<       鰑%@������������������������       �               ��/����?������������������������       �               E�JԮD!@�       �                 @���?����?       ��X�)B @������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?�       �                   �x�?�n��T�?       0~7�*@�       �                 �6Jy?�̥Q)�?       �9C�<�@�       �                 Њ�H?
4=�%�?       �(J��@�       �                    �?\n����?       � ��w<@������������������������       �               ��#���?�       �                 �j%?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               ��+��+@�       �                   s��?X�ߙ��?       /ʌu�h@�       �                 PK!�?�G���d�?        ��
��!G@�       �                 �C��?�L����?       Zk���>9@�       �                  Lm�?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?�       �                 �U��>��k���?       G+զm76@�       �                  �\�?d%@�"�?       ��[�@�       �                 ���?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               �cp>@������������������������       �        	       On��O0@�       �                 (I��?��^WJ�?       �=i�Z5@�       �                 0��?�[��Q��?       �\��#2@�       �                 zy?�?���_��?       x@���,(@�       �                 hU�<?H��aB��?       ����"@�       �                ��ߜ?L� P?)�?       ����x�@�       �                   .p�?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?������������������������       �               ��#�� @�       �                 P���?Ȕfm���?       ��Z�N@������������������������       �               ��#���?�       �                 0�C�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               H�4H�4@������������������������       �      �<       �cp>@�       �                 0��?�R{����?_       ����b@�       �                  `<��?����2��?$       f�vM@�       �                 `���?�5]���?       �ÖjD@�       �                 ��a?d�ߌv
�?       dXB@�       �                 �UaG?"7A ��?       r��¼�9@�       �                  ����?w>u���?       �+P7��2@�       �                 H��?,Lj����?       ���T�@������������������������       �               ;��,��@�       �                 Xnw�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?�       �                  ���?�� ��?       qp� k'@������������������������       �               0#0# @�       �                 ȯ�?���mf�?       毠�?b#@������������������������       �               �cp>@�       �                 0��?~�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @�       �                  ���?      �<       ���-��@������������������������       �               ��/����?������������������������       �               �cp>@�       �                 ���?�^�F�M�?	       ��ޚ�&@������������������������       �               ��+��+$@������������������������       �      ȼ       ��/����?�       �                 P3"!?      �<       ��#��@������������������������       �               ��#�� @������������������������       �               ��#�� @�       �                 ��?f/
�?       -���21@������������������������       �      �<       H�4H�4(@�       �                 �G��?     ��?       "F�b@������������������������       �               ��#�� @������������������������       �               H�4H�4@�       �                 p|߰?��z�Tf�?;       #aؕMW@�       �                 Џ��?�
^,��?       �鍅��<@�       �                 P��?j�4���?	       �.ex�^-@�       �                  �Mm�?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?�       �                 �`��?���mf�?       寠�?b#@������������������������       �      ��       ��/���@������������������������       �               0#0# @�       �                  ���?��p\�?       �����J,@������������������������       �               ��8��8*@������������������������       �      �<       ��#���?�       �                 �|'�?4��
|�?*       	��v\P@�       �                  ���?��'#�S�?       M��&GC@�       �                 �>J�?J����?       �N60@�       �                 pl8�?�'z�3�?
       ���da�%@�       �                 ��[M?h����?	       �����!@�       �                 `�[�?z��`p��?       �����@������������������������       �               H�4H�4@�       �                 `��?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?�       �                 �?�|2N��?       �3K}@������������������������       �               0#0# @������������������������       �               z�5��@�       �                   ���?���9�?       �q�Ί#6@�       �                @����?|��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �      ��       ��)��)3@������������������������       �               ��8��8:@�t�b�T     h�hhK ��h��R�(KK�KK��h �B8  �k(��b@hW�v%�f@aF`�a@���b:�^@����/k_@H�4H�48@��b:��Z@���|NV@H�4H�4@B����R@�H��tXU@H�4H�4@z�5��@�cp>7@        ;��,��@�cp>@        ��#�� @�cp>@        ��#�� @��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#���?                        ��/����?        z�5��@                ��#���?&jW�v%4@                'jW�v%4@        ��#���?                j1��tVQ@1����-O@H�4H�4@v�}wL@�+Q��B@0#0#�?]Lg1��F@��/���.@        \Lg1��&@���-��*@        �k(��"@�cp>@        z�5��@0����/@                0����/@        z�5��@                z�5��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ��#��@                ��#�� @��/���@        ��#���?                ��#���?��/���@                �cp>@        ��#���?��/����?        ��#���?                        ��/����?        Ey�5A@��/����?        �k(���5@                z�5��(@��/����?        \Lg1��&@                ��#���?��/����?                ��/����?        ��#���?                [Lg1��&@h
��6@0#0#�?��#���?��/���.@        ��#���?���-��@                ���-��@        ��#���?                        E�JԮD!@        ;��,��$@���-��@0#0#�?��#�� @���-��@0#0#�?        �cp>@0#0#�?        �cp>@                        0#0#�?��#�� @��/����?                ��/����?        ��#�� @                ��#�� @                z�5��(@��On�8@0#0# @z�5��@��/����?                ��/����?        z�5��@                z�5��@�e�_��7@0#0# @��#���?0����/3@        ��#���?                        /����/3@        ;��,��@0����/@0#0# @;��,��@0����/@                ��/����?        ;��,��@�cp>@                �cp>@        ;��,��@                                0#0# @���b:@@��/���@H�4H�4@z�5��8@                ���>��@��/���@H�4H�4@��#���?�cp>@0#0#�?��#���?                        �cp>@0#0#�?                0#0#�?        �cp>@        z�5��@��/����?0#0# @z�5��@        0#0#�?z�5��@                                0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?�P^Cy/@;l��F:B@vb'vb'2@��b:��*@�-����@@��+��+$@���>��@�]�ڕ�?@��+��+$@��#���?                z�5��@�]�ڕ�?@��+��+$@z�5��@鰑5@��+��+$@��#���?;l��F:2@0#0#@                0#0# @��#���?:l��F:2@0#0# @        D�JԮD1@0#0# @        ��/���@0#0# @        ��/����?0#0# @        ��/����?0#0#�?        ��/����?                        0#0#�?                0#0#�?        �cp>@                ���-��*@                D�JԮD!@                0����/@        ��#���?��/����?                ��/����?        ��#���?                ;��,��@�cp>@H�4H�4@                H�4H�4@;��,��@�cp>@H�4H�4@        �cp>@H�4H�4@        ��/����?                ��/����?H�4H�4@        ��/����?0#0#�?                0#0#�?        ��/����?                        0#0# @;��,��@                ��#���?                ��#��@                        鰑%@                ��/����?                E�JԮD!@        z�5��@��/����?        z�5��@                        ��/����?        ��#�� @�cp>@0#0# @��#�� @�cp>@H�4H�4@��#�� @�cp>@        ��#�� @��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                        ��/����?                        H�4H�4@                ��+��+@�#���9@�a#6�K@��~���\@�k(��"@���-��:@��+��+$@��#��@鰑5@        ��#�� @��/����?        ��#�� @                        ��/����?        ��#�� @'jW�v%4@        ��#�� @��/���@        ��#�� @��/����?                ��/����?        ��#�� @                        �cp>@                On��O0@        ;��,��@�cp>@��+��+$@;��,��@�cp>@��+��+$@;��,��@�cp>@0#0#@;��,��@�cp>@0#0#�?��#��@        0#0#�?��#�� @        0#0#�?��#�� @                                0#0#�?��#�� @                ��#���?�cp>@        ��#���?                        �cp>@                ��/����?                ��/����?                        H�4H�4@                H�4H�4@        �cp>@        ��#��0@��|��<@�o��oyZ@|�5��(@��/���.@�A�A>@<��,��$@��/���.@�A�A.@z�5��@��/���.@�A�A.@z�5��@��|��,@��+��+@z�5��@��/���@��+��+@z�5��@        0#0#�?;��,��@                ��#���?        0#0#�?��#���?                                0#0#�?        ��/���@0#0#@                0#0# @        ��/���@0#0# @        �cp>@                ��/����?0#0# @        ��/����?                        0#0# @        ���-��@                ��/����?                �cp>@                ��/����?��+��+$@                ��+��+$@        ��/����?        ��#��@                ��#�� @                ��#�� @                ��#�� @        �A�A.@                H�4H�4(@��#�� @        H�4H�4@��#�� @                                H�4H�4@��#��@���-��*@�i��R@��#���?D�JԮD!@��)��)3@        D�JԮD!@H�4H�4@        ��/����?0#0#@                0#0#@        ��/����?                ��/���@0#0# @        ��/���@                        0#0# @��#���?        ��8��8*@                ��8��8*@��#���?                z�5��@0����/@�C=�C=L@z�5��@0����/@�A�A>@z�5��@��/���@vb'vb'"@        ��/���@�C=�C=@        ��/����?�C=�C=@        ��/����?0#0#@                H�4H�4@        ��/����?0#0#�?        ��/����?                        0#0#�?                H�4H�4@        ��/����?        z�5��@        0#0# @                0#0# @z�5��@                        ��/����?��-��-5@        ��/����?0#0# @                0#0# @        ��/����?                        ��)��)3@                ��8��8:@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ:d�hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK兔h��B2         �                 0�0�?I�뎑.�?&      �A�>�~}@       �                 `��a?���;D��?�       �7`P�t@       �                 0�B�?�RY�w�?�       �/�s@       �                  K��?�W�/�h�?�       hE�]��p@       |                 ����?�b/ƃ:�?�       ��0k+p@                          �G�?��!�u�?�       ���2�m@                        0�X�?ny8�n�?       >l�~]G@                           �?��tV�?       �����B@	                        �sM?�#�8b�?       �Ǣ�98@
                        �?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?                        @߻V?      �<       %jW�v%4@������������������������       �               ��/����?������������������������       �        
       /����/3@                        ���>xf�T6|�?       y,*��P+@������������������������       �               ��#���?                        p���?�L����?       Yk���>)@������������������������       �               ��/���@                        赮�?
4=�%�?       �(J��@������������������������       �               ��#�� @������������������������       �               �cp>@                         ׃~?� �_rK�?       J�@��"@������������������������       �               z�5��@                        �N��?d%@�"�?       ��[�@������������������������       �      ��       ��/���@������������������������       �               ��#�� @       O                 �pur?n�ȿ��?m       ��4�h@       "                 �`>R?α��,��?B       D��[�^@       !                 �/��?Έ�-X�?	       q����2@                         �
;E?Ȕfm���?       ��Z�N/@������������������������       �               ��#��@������������������������       �               �cp>'@������������������������       �      ȼ       z�5��@#       :                    �?V�$�t�?9       gJ��Z@$       7                  �!�?� $hn�?)       ��oe"�S@%       (                   .p�?��9���?'       �o����R@&       '                 ��A?� �_rK�?       J�@��"@������������������������       �               ��/���@������������������������       �      ��       ;��,��@)       0                   ��?��#�ݬ?"       0X{Z�P@*       /                  ��d�?�N�'��?       �2WdK@+       .                 ��aӾ�hK)�?
       �h��K�2@,       -                  ����?�����?       �O��@������������������������       �      �<       ;��,��@������������������������       �      ȼ       ��/����?������������������������       �      �<       z�5��(@������������������������       �               �YLg1B@1       6                  ���?����X��?       &��֞&@2       3                `��0?`n����?       � ��w<@������������������������       �               ��#���?4       5                 ���Q?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#�� @8       9                p�	Y�?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?;       @                 0��{?��U�'�?       $��J��8@<       ?                 �΢뾌�6L�n�?       �E#��h @=       >                 8��p?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               z�5��@A       L                 �N�p?b��jʄ�?       @��m�0@B       I                 ����?ê��[�?	       @���`-@C       D                 �5W�?�̥Q)�?       �9C�<�@������������������������       �               �cp>@E       F                 0��>     ��?       "F�b@������������������������       �               0#0# @G       H                ���?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?J       K                �g ?      �<       ���-��@������������������������       �               ��/����?������������������������       �               0����/@M       N                  @mj�?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?P       k                 Ш��?���J�?+       �AJsQ@Q       T                   E(�?�w��?       �H�
�G@R       S                 ���2?��6L�n�?       �E#��h @������������������������       �      �<       ���>��@������������������������       �      ȼ       ��/����?U       h                 0S�r?��Iގ��?       �ܿtΠC@V       g                 g�a? ҿCB�?       �[�xA@W       Z                 �5�z?�R�u-��?       -=kD\=@X       Y                  �T?�����?       �O��@������������������������       �               ��/����?������������������������       �               ;��,��@[       f                  �j?8s���m�?       h[�ɝ97@\       e                 �{�?�m:�4�?       ���-X)@]       d                    �?l@ȱ��?       nm���S'@^       a                  �G?�?d%@�"�?       ��[�@_       `                 ��ߧ?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @b       c                 �e��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �      �<       鰑%@������������������������       �               0����/@i       j                 0��|?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?l       s                  �@�?�3O��?       s�W6@m       p                 P�M�?x���X��?
       (��֞&@n       o                 �~��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?q       r                 P�w?      �<       �k(��"@������������������������       �               ��#���?������������������������       �               ��#�� @t       u                  @?��?@b����?       �}IS&@������������������������       �               ;��,��@v       {                 ��h�?�� ��?       qp� k@w       z                 �v��?���mf�?       寠�?b@x       y                 �CK�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       �cp>@������������������������       �               0#0#�?}       �                      ��WT�V�?       D$_]3@~                           �?��6L�n�?	       �E#��h0@������������������������       �      �<       z�5��(@�       �                  �a�?���/��?       V��7�@������������������������       �               ��/����?�       �                 Z���?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?�       �                 �l�}?~%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 p��?H�F���?       :�.�-'@������������������������       �               鰑%@������������������������       �      �<       ��#���?�       �                 h��1?�K�"�^�?       �5
��wA@�       �                 ȯ�?�lRxN_�?       ��Ti�#>@������������������������       �               ��/����?�       �                 @Z˲?�I��'��?       ��u8<@�       �                 p�z�?��i���?       ����1@������������������������       �               ��+��+@�       �                 ����?Hy��]0�?	       ���y"(@������������������������       �               ��/����?�       �                  \��?�^�F�M�?       ��ޚ�&@������������������������       �               ��/����?������������������������       �               ��+��+$@�       �                 Q�?D5җ���?
       �E�=�X&@������������������������       �               z�5��@������������������������       �               0#0# @�       �                 Pր�?      �<       0����/@������������������������       �               ��/����?������������������������       �               �cp>@�       �                  `���?Ԛ�`p��?       T����=@�       �                 ��@�?���mf�?       毠�?b#@�       �                  �"�?�;[��G�?       �O�;�]!@�       �                 *�}?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                    �?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/���@������������������������       �               0#0#�?�       �                   +Y�?�?�0�!�?       a`�T�4@�       �                 ���?d����?       �����!@�       �                 0#ή?�v�;B��?       ՟���	 @�       �                    �?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?������������������������       �               #0#0&@�       �                 `�4x?�ޓ@���?Z       &��a@�       �                 P�f�?2�I�D��?+       ���[`Q@�       �                 ���?D}����?)       �J�j�P@�       �                   �x�?�djH�E�?       _�\m�n(@�       �                  �a�?�wV����?       Bi�i�"@������������������������       �               ��#�� @������������������������       �               0#0#�?�       �                 ��]?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?�       �                 Џ�B?J���d��?!       �co��J@�       �                 0�C�?�/E�
�?       �1��$7@�       �                 ����?��M�-�?
       �\�&�.@������������������������       �               ;��,��$@�       �                 @'��?hutee�?       Q9��@������������������������       �      �<       ��/����?������������������������       �               H�4H�4@�       �                 ���?���`�?       ��
�Me@�       �                   ��?��n��?       �-H�\@�       �                 ����?B��NV=�?       �t�ܲ@�       �                 @If�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                    �?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               0#0#�?�       �                 ��խ?`Da%��?       E���*=@�       �                 8�ۨ?m1�Q7�?       �5�T��%@�       �                 �I�W?<�a
=�?       ��l��@�       �                 �ԥ�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/���@������������������������       �               0#0#�?�       �                 p���?j,���O�?       ���/>@������������������������       �               H�4H�4@������������������������       �               ��#���?�       �                 �~��?H-����?
       hM��F2@������������������������       �               ��|��,@�       �                 ��K�?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �      �       ��+��+@�       �                 `���?(���?/       k!�#4�P@�       �                 p���?�,�c���?*       �Km X;N@�       �                 PiU�?d*�'=P�?        �2"@������������������������       �               0#0# @������������������������       �      ȼ       ��/����?������������������������       �      ��#       ~˷|˷I@�       �                 H��?�AP�9��?       i��6��@������������������������       �               H�4H�4@�       �                 @���?|�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @�t�bh�hhK ��h��R�(KK�KK��h �Bx  �k(���e@`�ڕ��d@?��8�c`@g:��,&c@	���|�`@[��Y��H@g:��,&c@��/���^@�s?�s?=@1�����b@��h�\@H�4H�4@�k(��b@�cp>�Y@H�4H�4@�5�װ`@��On�X@H�4H�4@�k(��"@�+Q��B@        ��#��@�-����@@        ��#���?�cp>7@        ��#���?�cp>@                �cp>@        ��#���?                        %jW�v%4@                ��/����?                /����/3@        z�5��@鰑%@        ��#���?                ��#�� @鰑%@                ��/���@        ��#�� @�cp>@        ��#�� @                        �cp>@        ;��,��@��/���@        z�5��@                ��#�� @��/���@                ��/���@        ��#�� @                �P^Cy_@3����-O@H�4H�4@:��P^�V@�_��e�=@H�4H�4@���>��@�cp>'@        ��#��@�cp>'@        ��#��@                        �cp>'@        z�5��@                >��,��T@:l��F:2@H�4H�4@������Q@��/���@        j1��tVQ@�cp>@        ;��,��@��/���@                ��/���@        ;��,��@                ���b:P@��/����?        ��b:��J@��/����?        ��,���1@��/����?        ;��,��@��/����?        ;��,��@                        ��/����?        z�5��(@                �YLg1B@                ;��,��$@��/����?        ��#�� @��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                ��#�� @                ��#�� @��/����?        ��#�� @                        ��/����?        [Lg1��&@鰑%@H�4H�4@���>��@��/����?        ��#���?��/����?                ��/����?        ��#���?                z�5��@                ��#��@0����/#@H�4H�4@��#�� @0����/#@H�4H�4@��#�� @�cp>@H�4H�4@        �cp>@        ��#�� @        H�4H�4@                0#0# @��#�� @        0#0#�?��#�� @                                0#0#�?        ���-��@                ��/����?                0����/@        ��#�� @                ��#���?                ��#���?                Fy�5A@Pn��O@@H�4H�4@�k(��2@�a#6�;@0#0#�?���>��@��/����?        ���>��@                        ��/����?        [Lg1��&@���-��:@0#0#�?���>��@�cp>�9@0#0#�?���>��@鰑5@0#0#�?;��,��@��/����?                ��/����?        ;��,��@                ��#�� @%jW�v%4@0#0#�?��#�� @0����/#@0#0#�?��#�� @/����/#@        ��#�� @��/���@        ��#�� @��/����?                ��/����?        ��#�� @                        �cp>@                ��/����?                ��/����?                �cp>@                        0#0#�?        鰑%@                0����/@        ��#��@��/����?        ��#��@                        ��/����?        �P^Cy/@0����/@0#0# @<��,��$@��/����?        ��#���?��/����?                ��/����?        ��#���?                �k(��"@                ��#���?                ��#�� @                ;��,��@��/���@0#0# @;��,��@                        ��/���@0#0# @        ��/���@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@                        0#0#�?�P^Cy/@��/���@        ���>��,@��/����?        z�5��(@                ��#�� @��/����?                ��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#���?鰑%@                鰑%@        ��#���?                z�5��@D�JԮD!@%S2%S27@z�5��@��/���@%S2%S27@        ��/����?        z�5��@��/����?%S2%S27@        ��/����?�A�A.@                ��+��+@        ��/����?��+��+$@        ��/����?                ��/����?��+��+$@        ��/����?                        ��+��+$@z�5��@        0#0# @z�5��@                                0#0# @        0����/@                ��/����?                �cp>@                0����/#@��+��+4@        ��/���@0#0# @        ��/���@0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                �cp>@                ��/����?                ��/���@                        0#0#�?        ��/����?vb'vb'2@        ��/����?�C=�C=@        ��/����?�C=�C=@        ��/����?0#0#�?                0#0#�?        ��/����?                        H�4H�4@        ��/����?                        #0#0&@<��,��4@E�JԮDA@�N��NlT@<��,��4@�]�ڕ�?@S2%S2%1@<��,��4@�]�ڕ�?@H�4H�4(@��#�� @��/����?0#0# @��#�� @        0#0#�?��#�� @                                0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?|�5��(@�_��e�=@��+��+$@\Lg1��&@���-��@��+��+@<��,��$@��/����?H�4H�4@;��,��$@                        ��/����?H�4H�4@        ��/����?                        H�4H�4@��#���?0����/@0#0# @��#���?0����/@0#0#�?��#���?��/����?0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?��#���?��/����?                ��/����?        ��#���?                        �cp>@                        0#0#�?��#���?�cp>7@��+��+@��#���?�cp>@0#0#@        �cp>@0#0#�?        �cp>@                ��/����?                ��/���@                        0#0#�?��#���?        H�4H�4@                H�4H�4@��#���?                        E�JԮD1@0#0#�?        ��|��,@                �cp>@0#0#�?                0#0#�?        �cp>@                        ��+��+@        �cp>@2#0#P@        ��/����?����M@        ��/����?0#0# @                0#0# @        ��/����?                        ~˷|˷I@        ��/����?��+��+@                H�4H�4@        ��/����?0#0# @        ��/����?                        0#0# @�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�I]fhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKㅔh��B�1         �                 ���b?.�O��N�?-      -�mLc�}@       �                  �l�?ef�����?�       OY�,K<u@       �                 �
o?߬��a�?�       C�v�[t@       u                 ��^�?%k��?�       ����	l@       4                 h�"d?P�����?~       �)�$�&h@       #                 ��?�\#�C�??       0`R;Z@                          \��?�HU����?       "��N��E@                        �T�
?���(x�?       �B�n:@	       
                 `���>`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#��@                        �2�Y?�`@s'��?       �[�_4@                           �?f%@�"�?       ��[�@                        P@t.?& k�Lj�?       �q��l}@������������������������       �               �cp>@                        *#�g?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#���?                        ���R?��&���?       ��G2��,@������������������������       �               ���-��*@������������������������       �      �<       ��#���?                         �b'�?r����?       $c�Z%K1@                        8T��?M�����?       p����.@                        �y�����=�Sο?
       ����,@                        ���>`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?                         ��d�?      �<       [Lg1��&@������������������������       �               ��#�� @������������������������       �               �k(��"@������������������������       �      ȼ       ��/����?!       "                  P�"�?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?$       1                 @*tC?�d�$���?"       ?��#�N@%       0                 �؉�?�LI)Z��?       Ji_y,*K@&       /                   ��?�,AF@��?       ^k���>I@'       .                  �~��? u.?��?       Ω��`�:@(       +                  W�5?���P��?       �*Y�ȹ9@)       *                 �r��?�q�Ptܳ?       P�� 5�7@������������������������       �      ȼ       \Lg1��6@������������������������       �      �<       ��/����?,       -                    �?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               �,����7@������������������������       �      ȼ       ��/���@2       3                 ��f�?��|��?       ���ĺw@������������������������       �               0����/@������������������������       �               ��#�� @5       <                 ���?����_�??       V�_9�V@6       7                 �/��?�^�#΀�?       P�{��A5@������������������������       �               ��#���?8       9                 �j%?��٤ݸ?
       ��<5�84@������������������������       �               ���-��*@:       ;                 PeT�?�`@s'��?       Ei_y,*@������������������������       �               �cp>@������������������������       �               ��#���?=       b                 �U��>`��jʄ�?4       A��m�P@>       K                 �!�?�A���?       ,J�7��?@?       J                 @�Ǻ?憛���?	       �7vg�#@@       A                 �v�(?���`�?       ��
�Me@������������������������       �               ��#���?B       I                 �ҭ?��[����?       Il�_A@C       H                 �~�?~�G���?       ��%�|@D       E                 �X��?|��`p��?       �����@������������������������       �               0#0#�?F       G                 �u+�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               �cp>@������������������������       �               0#0# @L       Y                 0C�?_9D��?       C.�|6@M       R                 ��-�?\n����?       Ԁh��K.@N       Q                  P���?$ k�Lj�?       �q��l}@O       P                 ���Y?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               �cp>@S       V                   \��?�FO���?       �ߌ$@T       U                 `ಣ?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ���>��@W       X                 ��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?Z       _                 ���?��d
���?       f�G�N�@[       ^                 �j�?����|e�?       �z �B�@\       ]                 �Z�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0# @`       a                 ����?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?c       l                 0��?ԢV���?       mk;{�A@d       g                 P
��?�8f���?       ֑+XW�+@e       f                 �j�Y?X�r{��?       e�6� @������������������������       �               ���-��@������������������������       �               ��#���?h       k                 n�
Q?Hy��]0�?       ���y"@i       j                 p��?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0#@m       n                 �ĕ�?X�+���?       �aJ9U5@������������������������       �               ��#���?o       r                  P���?�3+�Pr�?       [-"�=L4@p       q                 �=��?      �<	       ��On�(@������������������������       �               �cp>@������������������������       �               /����/#@s       t                 ��A�?��fm���?       ��Z�N@������������������������       �               ��#�� @������������������������       �               �cp>@v       w                 P8��?v�p�?       ����>?@������������������������       �               H�4H�4(@x       �                 H���?tL�0���?       Q~�)��2@y       z                   .p�?֘�?ʊ�?	       ��l���)@������������������������       �               �cp>@{       �                 @Z˲?ھ�R���?       :�S) $@|       }                  t�?X*�'=P�?        �2"@������������������������       �               H�4H�4@~                        �fQ?z��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �      �<       ��#���?������������������������       �               H�4H�4@�       �                  	͖?�q��?A       ����lXY@�       �                 ���?H�I���?'       G*��Z�O@�       �                 ��I�? �W�W��?       �Zc���8@�       �                 ��~?꜋���?       aJ9U63@�       �                  ;��?2�c3���?       �uk��!@������������������������       �               �cp>@�       �                 ��J?^n����?       � ��w<@�       �                 T�@?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �               z�5��@�       �                 ����?�FO���?       �ߌ$@������������������������       �      �<       ���>��@�       �                 X���?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      �<       �cp>@�       �                      d))5���?       �|�xhcC@�       �                  `���?�Lh� ��?       Ƚ�@��?@������������������������       �               �k(���5@�       �                 �Mr�?
����?       ���"�X$@������������������������       �      �<       ���>��@�       �                 �~�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                  `�J�?��|��?       ���ĺw@������������������������       �               0����/@������������������������       �               ��#�� @�       �                 �*��?���\z_�?       ��e~�B@�       �                 ��?إ�je��?       ��BLGh0@�       �                 0��?h�4���?       �tCP��@������������������������       �               0#0# @������������������������       �               �cp>@������������������������       �               �cp>'@�       �                 `(¢?�Z�����?       U�N�:5@�       �                  �[??x�����?	       �iO9T�.@�       �                  ���?l����?       P	K��,@������������������������       �               ��/����?�       �                 ��y�?`�s�	�?       e���*@������������������������       �      ��       z�5��(@������������������������       �      ȼ       ��/����?������������������������       �               0#0#�?�       �                 @mo�?��íxq�?       $2��-�@�       �                 �C8�?�@G���?       hu��@�       �                  R��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 ���H?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 �\��?��!��?       �@��&,@�       �                 (�*�?�/y߃�?
       Ɓ\��((@������������������������       �               ��#���?�       �                 �:WN?�^�F�M�?	       ��ޚ�&@������������������������       �               0#0# @�       �                 ��
�?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 ��ǩ?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                    �?�_$��g�?P       �7�?0�`@�       �                  p<��?H,�}��?%       ��2P4L@������������������������       �               ��#���?�       �                 �å�?8>�fn �?$       �z���K@�       �                   E(�?�n���k�?       3��&�:@�       �                  f!�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               %S2%S27@������������������������       �      �<       �s?�s?=@�       �                 �p^�?�k��*��?+       2�p�W�R@�       �                 0��?��[����?       Hl�_A@������������������������       �               0#0#�?�       �                 p�҇?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �               0����/@�       �                 @�?@͈+���?'       l��AFQ@�       �                 ����?<4�}���?&       �C�u�P@�       �                 ���?��H�&p�?       N^�3��E@������������������������       �        	       0#0#0@�       �                 pL�s?�AP�9��?       i��6��;@������������������������       �               ��/���@�       �                 `%�?Ny��]0�?       ���y"8@�       �                 �-�?�T`�[k�?
       �m����0@�       �                 p�Z�?��E�B��?	       dߞKC.@�       �                 ���?t��ճC�?       y��l$,@�       �                 p��?|��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               #0#0&@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?������������������������       �               �C=�C=@������������������������       �               %S2%S27@������������������������       �      �<       ��/����?�t�bh�hhK ��h��R�(KK�KK��h �BH  C����b@O��+c@׬�ڬe@1�����b@��t�Ha@������J@�#���b@�-����`@�
��
�E@;��P^�V@�e�_��W@��)��)C@�GpAV@�cp>W@H�4H�4(@��,���Q@F�JԮDA@        <��,��4@�cp>7@        ���>��@0����/3@        ��#��@��/����?                ��/����?        ��#��@                z�5��@D�JԮD1@        ��#�� @��/���@        ��#���?��/���@                �cp>@        ��#���?��/����?        ��#���?                        ��/����?        ��#���?                ��#���?���-��*@                ���-��*@        ��#���?                ��b:��*@��/���@        ��b:��*@��/����?        ��b:��*@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        [Lg1��&@                ��#�� @                �k(��"@                        ��/����?                ��/����?                ��/����?                ��/����?        }�5��H@�cp>'@        �,����G@���-��@        �,����G@�cp>@        �,����7@�cp>@        �,����7@��/����?        \Lg1��6@��/����?        \Lg1��6@                        ��/����?        ��#���?��/����?                ��/����?        ��#���?                        ��/����?        �,����7@                        ��/���@        ��#�� @0����/@                0����/@        ��#�� @                �k(��2@��|��L@H�4H�4(@��#�� @0����/3@        ��#���?                ��#���?/����/3@                ���-��*@        ��#���?�cp>@                �cp>@        ��#���?                ��#��0@2����/C@H�4H�4(@|�5��(@��On�(@�C=�C=@��#���?0����/@0#0#@��#���?0����/@0#0# @��#���?                        0����/@0#0# @        ��/����?0#0# @        ��/����?0#0# @                0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?                �cp>@                        0#0# @\Lg1��&@��/���@H�4H�4@<��,��$@0����/@        ��#���?��/���@        ��#���?��/����?                ��/����?        ��#���?                        �cp>@        �k(��"@��/����?        ��#�� @                ��#���?                ���>��@                ��#���?��/����?        ��#���?                        ��/����?        ��#���?�cp>@H�4H�4@        ��/����?H�4H�4@        ��/����?0#0#�?                0#0#�?        ��/����?                        0#0# @��#���?��/����?                ��/����?        ��#���?                ��#��@�cp>�9@��+��+@��#���?��/���@��+��+@��#���?���-��@                ���-��@        ��#���?                        ��/����?��+��+@        ��/����?0#0#�?                0#0#�?        ��/����?                        0#0#@z�5��@:l��F:2@        ��#���?                ��#�� @:l��F:2@                ��On�(@                �cp>@                /����/#@        ��#�� @�cp>@        ��#�� @                        �cp>@        ��#���?��/���@��8��8:@                H�4H�4(@��#���?��/���@�C=�C=,@��#���?��/���@0#0# @        �cp>@        ��#���?��/����?0#0# @        ��/����?0#0# @                H�4H�4@        ��/����?0#0# @                0#0# @        ��/����?        ��#���?                                H�4H�4@���>��L@2����/C@��+��+@�GpAF@;l��F:2@0#0#�?��b:��*@�cp>'@        ��b:��*@�cp>@        ��#��@0����/@                �cp>@        ��#��@��/����?        ��#���?��/����?                ��/����?        ��#���?                z�5��@                �k(��"@��/����?        ���>��@                ��#�� @��/����?        ��#�� @                        ��/����?                �cp>@        �P^Cy?@���-��@0#0#�?���>��<@��/����?0#0#�?�k(���5@                ���>��@��/����?0#0#�?���>��@                        ��/����?0#0#�?                0#0#�?        ��/����?        ��#�� @0����/@                0����/@        ��#�� @                ��b:��*@%jW�v%4@0#0#@        ��|��,@0#0# @        �cp>@0#0# @                0#0# @        �cp>@                �cp>'@        ��b:��*@�cp>@0#0# @z�5��(@��/����?0#0#�?z�5��(@��/����?                ��/����?        {�5��(@��/����?        z�5��(@                        ��/����?                        0#0#�?��#���?��/���@0#0#�?        �cp>@0#0#�?        �cp>@                ��/����?                ��/����?                        0#0#�?��#���?��/����?        ��#���?                        ��/����?        ��#�� @��/����?��+��+$@��#���?��/����?��+��+$@��#���?                        ��/����?��+��+$@                0#0# @        ��/����?0#0# @        ��/����?                        0#0# @��#���?��/����?        ��#���?                        ��/����?        ��#���?On��O0@�[��[�\@��#���?��/����?������J@��#���?                        ��/����?������J@        ��/����?H�4H�48@        ��/����?0#0#�?                0#0#�?        ��/����?                        %S2%S27@                �s?�s?=@        ��|��,@.��+��N@        0����/@0#0# @                0#0#�?        0����/@0#0#�?                0#0#�?        0����/@                0����/#@����M@        ��/���@
����M@        ��/���@xb'vb'B@                0#0#0@        ��/���@��+��+4@        ��/���@                ��/���@��+��+4@        ��/���@��8��8*@        ��/����?��8��8*@        ��/����?��8��8*@        ��/����?0#0# @                0#0# @        ��/����?                        #0#0&@        ��/����?                ��/����?                        �C=�C=@                %S2%S27@        ��/����?        �t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�޵#hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKυ�h��BH-         x                 ��q�?F"���O�?%      #����u}@       s                 ���?b�j����?�       �g;�6q@       r                 �{?r�'%��?�       ���9�Tp@       Y                 P�}A?��g�r��?�        �6D�n@       N                    �?�(�؇��?z       �� уg@       +                  ��i?M���Ю�?e       ~�ޟ��c@                         �C
T?��bxv�?6       r'�3	lW@                        �C[?�^����?$       �Yk���O@	       
                  �{��?`�r{��?       e�6� /@������������������������       �      ��       ���-��*@������������������������       �               ��#�� @                        p��?fn����?       � ��w<H@                        ~`���̅����?       O� ���D@                        �"c?
��I@�?       �2d�%@                         /�`?X�r{��?       e�6� @������������������������       �               ��#���?                        (�!�?      �<       ���-��@������������������������       �               ��/����?������������������������       �               0����/@                        ��x?hn����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?                           �?�	�� ��?       @�x��>@������������������������       �               z�5��8@                        � �}?�����?       �O��@                        ĵ��>      �<       ��#��@������������������������       �               ��#�� @������������������������       �               ��#�� @                        0z��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      Լ       ���-��@!       "                  �Ԧ�?�N,u��?       ��u�=@������������������������       �               ��/����?#       (                 ���X?8Bms�?       ��֖��;@$       %                 ���?���OT�?       r�>%,�9@������������������������       �        
       ������3@&       '                 �?�����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?)       *                 @�C�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?,       3                 ����?�ٙJ���?/       �'%)P@-       .                 �_�?<3#܅�?       ���A�0@������������������������       �               ��#���?/       0                  @?��?`�r{��?       e�6� /@������������������������       �      м       D�JԮD!@1       2                 ��~?��|��?       ���ĺw@������������������������       �      ��       0����/@������������������������       �               ��#�� @4       5                 �N�p?\0�D���?"       ��yIgH@������������������������       �               ��+��+@6       K                 0
��?�tU��a�?        0���E@7       H                  �j?q����?       ؔn�vC@8       E                 ��d?�>dCQ�?       ��9ƞP;@9       D                  �G?�?4�Cx@��?       X�k�30@:       ;                 x��?ެͅV�?	       c�U(@������������������������       �               ��#�� @<       C                   ��?B�pB}��?       ����1$@=       B                   ���?��r�g��?       ��1ֻ�@>       A                   .p�?
4=�%�?       �(J��@?       @                 ���?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��#��@������������������������       �      м       ��/���@F       G                 �m۶?����X��?	       '��֞&@������������������������       �               ��/����?������������������������       �      �<       <��,��$@I       J                 q� ?h�ђ���?       �oFݜh%@������������������������       �               ��#�� @������������������������       �               D�JԮD!@L       M                    �?      �<       ��+��+@������������������������       �               0#0# @������������������������       �               H�4H�4@O       P                @0W=e?8�q�W�?       ~KoS�=@������������������������       �               ��/����?Q       X                 ����?�=�Sο?       ����<@R       S                  `���?�-�r?�?       �M�)#�;@������������������������       �               �,����7@T       U                 �Mr�?�����?       ��X�)B@������������������������       �               ��#�� @V       W                    �?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      �<       ��/����?Z       i                 ���O?C���(�?        � l�̅M@[       ^                 `�ռ?�O-r��?       �bY�RC@\       ]                 P>-l?@r�]i��?       ��U�i�9@������������������������       �               ��On�8@������������������������       �      �<       ��#���?_       `                @�-b!?`n����?       � ��w<(@������������������������       �               ��/����?a       b                 X��?���Ѯ�?       ��GQ&@������������������������       �               ;��,��@c       d                �s�ar?���/��?       @z$S��@������������������������       �               ��#�� @e       h                 ����?Ȕfm���?       ��Z�N@f       g                  @?��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��#���?j       q                   B�?邞ñ`�?       �;%��4@k       p                 h'v�?���Ul��?	        {|3�0@l       o                 �n6�?Ĕfm���?       �0��z'@m       n                 H�a�?��Z�	7�?       j~���@������������������������       �               z�5��@������������������������       �      �<       ��/����?������������������������       �      ��       ���-��@������������������������       �      �<       ;��,��@������������������������       �               0#0#@������������������������       �     ��
       �C=�C=,@t       u                  �Os?h�p\�?       �����J,@������������������������       �               ��+��+$@v       w                 v�?f,���O�?       ���/>@������������������������       �               H�4H�4@������������������������       �               ��#���?y       �                  �\�?����I�?{       �8���}h@z       �                 �7�?��%U�?       ,��q`i8@{       ~                 @tܣ?N^�GH�?       >cmiW6@|       }                  p�{�?��Z�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@       �                 -��?�0�~��?	       r��GQ1@������������������������       �               0#0#�?������������������������       �               On��O0@������������������������       �      �<       ��#�� @�       �                 ���? �,��?n       ����pe@�       �                  �Ԧ�?~��w��?0       ʠ3u�DR@�       �                  s�}?*���x��?       ����@@�       �                  MѴ?���uȇ�?       ��&"�8@������������������������       �               0#0#@�       �                 ����? ��x	��?       ��a�4@�       �                 �3�?�T�"��?       ��`2�Z+@������������������������       �               H�4H�4@�       �                 �_�?��XnP��?       ЭS`oM%@�       �                 P��?x5JH���?       �MOI#@�       �                 �Ċ?���mf�?       毠�?b@������������������������       �      �<       ��/���@������������������������       �               0#0#�?������������������������       �               0����/@������������������������       �               0#0#�?�       �                 �o|Q?�_�A�?       肵�e`@������������������������       �      �<       ;��,��@������������������������       �      ȼ       ��/����?������������������������       �               vb'vb'"@�       �                 ��0�?���~��?       �$JE��C@�       �                 pN�u?ڦ$Rď�?       �;h&:=@�       �                 ��:�?�3+�Pr�?       Z-"�=L4@�       �                 G҈n?      �<       0����/#@������������������������       �               ��/����?������������������������       �               ��/���@�       �                 pa��?R�ђ���?       �oFݜh%@������������������������       �               ��#�� @�       �                 0���?      �<       D�JԮD!@������������������������       �               �cp>@������������������������       �               �cp>@�       �                  `s�?z��`p��?       f;3@��!@������������������������       �               �cp>@������������������������       �      �<       H�4H�4@�       �                ��5p�?��AH�.�?       ���D��#@�       �                 ��?��d
���?       f�G�N�@�       �                 H�z�?����]L�?       N66�ͯ@�       �                 �m��?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               0#0# @������������������������       �               H�4H�4@�       �                 @�	�?��Sg��?>       ڐ�7�X@�       �                 �ʨ�?J�'��u�?'       u��>"�O@�       �                 �	I�?��i�#%�?#       �� �^�L@�       �                  �9��?ԉ:�j��?       �2Z�D@������������������������       �               ��#���?�       �                  ;��?��Z"�b�?       ]��Q�(D@������������������������       �               S2%S2%1@�       �                  ���?����	��?       eR�P�,7@�       �                    �?�~���9�?       �q�Ί#6@�       �                 �sh�?Hy��]0�?       ���y"@�       �                 �5Ry?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      ��       H�4H�4@������������������������       �               0#0#0@������������������������       �      �<       ��#���?�       �                  P�"�?|�h����?
       ��[�/@������������������������       �               ��/����?�       �                 �ˮ�?�j.�d��?	       �I���+@������������������������       �               ��+��+$@�       �                  ��?�@G���?       hu��@������������������������       �               ��/����?�       �                 @�C�?~�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 �U��?��q�R�?       C}Ԥ@�       �                 �{��?|�G���?       ��%�|@������������������������       �      �<       ��/����?������������������������       �               0#0# @������������������������       �               ��#�� @�       �                 ��?X�M��b�?       8��0��A@������������������������       �               �s?�s?=@�       �                 P�k�?���`p��?       �����@������������������������       �               ��/����?������������������������       �      ��       0#0#@�t�bh�hhK ��h��R�(KK�KK��h �Bh  �#���b@�)�B�d@��
���c@�P^CyM`@%�B��Y@��-��-E@�t�Y,`@&�B��Y@�s?�s?=@�t�Y,`@&�B��Y@�A�A.@.�����[@Pn��OP@#0#0&@���#8U@3����-O@#0#0&@��>���N@Pn��O@@        ��,���A@��|��<@        ��#�� @���-��*@                ���-��*@        ��#�� @                ��#��@@��/���.@        ��#��@@E�JԮD!@        z�5��@��/���@        ��#���?���-��@        ��#���?                        ���-��@                ��/����?                0����/@        ��#�� @��/����?        ��#�� @                        ��/����?        Jp�}>@��/����?        z�5��8@                ;��,��@��/����?        ��#��@                ��#�� @                ��#�� @                ��#���?��/����?                ��/����?        ��#���?                        ���-��@        �#���9@��/���@                ��/����?        
�#���9@��/����?        |�5��8@��/����?        ������3@                ;��,��@��/����?        ;��,��@                        ��/����?        ��#���?��/����?                ��/����?        ��#���?                �,����7@�_��e�=@#0#0&@z�5��@���-��*@        ��#���?                ��#�� @���-��*@                D�JԮD!@        ��#�� @0����/@                0����/@        ��#�� @                <��,��4@On��O0@#0#0&@                ��+��+@<��,��4@Nn��O0@H�4H�4@<��,��4@On��O0@0#0#�?�k(��2@��/���@0#0#�?��#�� @���-��@0#0#�?��#�� @�cp>@0#0#�?��#�� @                z�5��@�cp>@0#0#�?��#�� @�cp>@0#0#�?��#�� @�cp>@        ��#�� @��/����?        ��#�� @                        ��/����?                ��/����?                        0#0#�?��#��@                        ��/���@        ;��,��$@��/����?                ��/����?        <��,��$@                ��#�� @D�JԮD!@        ��#�� @                        D�JԮD!@                        ��+��+@                0#0# @                H�4H�4@��b:��:@�cp>@                ��/����?        ��b:��:@��/����?        ��b:��:@��/����?        �,����7@                z�5��@��/����?        ��#�� @                ��#���?��/����?                ��/����?        ��#���?                        ��/����?        ��,���1@�+Q��B@0#0#@�k(��"@��|��<@        ��#���?��On�8@                ��On�8@        ��#���?                ��#�� @��/���@                ��/����?        ��#�� @�cp>@        ;��,��@                z�5��@�cp>@        ��#�� @                ��#���?�cp>@                �cp>@                ��/����?                ��/����?        ��#���?                ��#�� @E�JԮD!@0#0#@��#�� @D�JԮD!@        z�5��@E�JԮD!@        z�5��@��/����?        z�5��@                        ��/����?                ���-��@        ;��,��@                                0#0#@                �C=�C=,@��#���?        ��8��8*@                ��+��+$@��#���?        H�4H�4@                H�4H�4@��#���?                ��,���1@1����-O@��~���\@;��,��@:l��F:2@0#0#�?z�5��@:l��F:2@0#0#�?z�5��@��/����?                ��/����?        z�5��@                        On��O0@0#0#�?                0#0#�?        On��O0@        ��#�� @                z�5��(@h
��F@�[��[�\@��#�� @E�JԮDA@�A�A>@;��,��@鰑%@vb'vb'2@;��,��@鰑%@vb'vb'"@                0#0#@;��,��@鰑%@��+��+@        E�JԮD!@��+��+@                H�4H�4@        E�JԮD!@0#0# @        D�JԮD!@0#0#�?        ��/���@0#0#�?        ��/���@                        0#0#�?        0����/@                        0#0#�?;��,��@��/����?        ;��,��@                        ��/����?                        vb'vb'"@z�5��@�e�_��7@H�4H�4(@��#�� @鰑5@H�4H�4@��#�� @:l��F:2@                0����/#@                ��/����?                ��/���@        ��#�� @D�JԮD!@        ��#�� @                        D�JԮD!@                �cp>@                �cp>@                �cp>@H�4H�4@        �cp>@                        H�4H�4@��#���?�cp>@H�4H�4@��#���?�cp>@H�4H�4@��#���?�cp>@0#0#�?��#���?        0#0#�?                0#0#�?��#���?                        �cp>@                        0#0# @                H�4H�4@��#��@/����/#@��-��-U@��#��@��/���@�˷|˷I@��#�� @�cp>@\��Y��H@��#�� @��/����?��)��)C@��#���?                ��#���?��/����?��)��)C@                S2%S2%1@��#���?��/����?��-��-5@        ��/����?��-��-5@        ��/����?��+��+@        ��/����?0#0# @        ��/����?                        0#0# @                H�4H�4@                0#0#0@��#���?                        0����/@#0#0&@        ��/����?                �cp>@#0#0&@                ��+��+$@        �cp>@0#0#�?        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?��#�� @��/����?0#0# @        ��/����?0#0# @        ��/����?                        0#0# @��#�� @                        ��/����?B�A�@@                �s?�s?=@        ��/����?0#0#@        ��/����?                        0#0#@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�G�hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK兔h��B2         f                 0C�?�qaWF�?#      ��r��}@       O                 ��??�-K��>�?�       ��@��>m@       6                 `8s�?�IɁ�-�?h       ]E���f@       #                 �U���jF>(���?G       �EBCZH^@                           �?�-����?!       ^�:&L@                          ��?�3���r�?       X�i�ҺC@������������������������       �               ��/���@                          p��?vU�vѢ�?       lӶ��A@	       
                  �JV�?V�'r��?       �
$�TA@������������������������       �               �k(��"@                        ��w?lzw��?       �B޳�X9@                        ���d?   ���?	       *x�1�)@                         Pmj�?Zn����?       ~��Y-"@������������������������       �               ��/����?                        x��?T����?       Q	K��@������������������������       �      �<       ;��,��@                        ��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      м       ��/���@������������������������       �      ��       z�5��(@������������������������       �      �<       ��/����?                         �)�?�z���`�?       �7���0@                        ��t?�PJo�x�?       V|qt�&@                         8hV?& k�Lj�?       �q��l}@������������������������       �               ��/����?                        �$I�?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?                        ����?�����?       �O��@������������������������       �               ��/����?������������������������       �      �<       ;��,��@!       "                 @Ws�?t@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@$       %                 ���#?�Gk���?&       ٖ��<5P@������������������������       �               Dy�5A@&       1                 �p�?�����?       �h�d��>@'       .                  �x��?h�s�	�?       h���:@(       -                 �N4m?\����?       P	K��,@)       ,                 �~�?�_�A�?       炵�e`@*       +                 �L'?�����?       �O��@������������������������       �               ��/����?������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?������������������������       �               ���>��@/       0                  1�>      �<	       |�5��(@������������������������       �               ��#���?������������������������       �               [Lg1��&@2       3                  �~��?ޔfm���?       ��Z�N@������������������������       �               ��/����?4       5                    �?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?7       @                  ㌇?�x�x��?!       �����K@8       9                 �V��?Ȕfm���?       3�x�А3@������������������������       �               /����/#@:       =                �3�.s?���/��?       6��o��#@;       <                 P�f�?, k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      �<       ��/���@>       ?                 T��p?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@A       H                 �_��?u#N��?        �b�"B@B       G                  ��d�?z�G���?	       '5L�`�'@C       D                 �m۶?�;�a
=�?       ��l��@������������������������       �               0����/@E       F                  �j?z�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               ��+��+@I       N                 �O��?��x_F-�?       x%jW�v8@J       K                 D��?�:�^���?       ��]�ڕ5@������������������������       �               ��#��0@L       M                 `iY�?�Z�	7�?       i~���@������������������������       �      ȼ       ��/����?������������������������       �               z�5��@������������������������       �      �<       �cp>@P       c                 hJ��?TO{��A�?&       ���v8L@Q       ^                  7u�?�_�ѡ��?       �`��|H@R       [                 �l�}?d�4��d�?       ,�V��vC@S       V                 @F�.>櫐�?       ��j���6@T       U                 �S�?��Tu��?       ����.@������������������������       �      ��
       ��|��,@������������������������       �      ܼ       ��#���?W       Z                 8��?�_�A�?       肵�e`@X       Y                    �?�����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?\       ]                 �%N�?إ�je��?       ��BLGh0@������������������������       �      ��       ��|��,@������������������������       �               0#0# @_       `                 0eŎ?�Z�	7�?       j~���$@������������������������       �               ;��,��@a       b                 �L�I?& k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      �<       ��/���@d       e                 �	��?�w�;B��?       ՟���	 @������������������������       �               �C=�C=@������������������������       �      ȼ       ��/����?g       �                   ��?������?�       /��:I�m@h       �                 0���?-C]��?e       �-�
ld@i       r                 �N�p?�yh���?&       ��>\1O@j       k                   ��?a{���?       �~8�31@������������������������       �               ��/����?l       q                 pM�?$ȇ��?       ��8.@m       p                 �ˌ}?�K��t�?       M����"@n       o                    �?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0#@������������������������       �               z�5��@������������������������       �               H�4H�4@s       ~                 NK�X?��Bt{�?       R�"���F@t       u                 ��f�?�Wf]�?       ?���g�!@������������������������       �               ��#���?v       }                 p>r�?�~�&��?       @�]��@w       |                 0J(�?l�4���?       �tCP��@x       y                 �U�,?�@G���?       hu��@������������������������       �               0#0#�?z       {                    �?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               H�4H�4@       �                  ���?.���?       @�w�&3B@������������������������       �               ��/���@�       �                 ����?b�p����?       T�Ĭ�G@@�       �                 �F�{?U�}R4�?       �[RZ��#@������������������������       �               ��#�� @�       �                 0&�r?�1�RH3�?       <�����@�       �                 p� �?��íxq�?       $2��-�@�       �                  �P�?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �      ��       ��/���@������������������������       �               0#0# @�       �                 �^J�? ��'��?       ��_�
�6@�       �                 pTF�?�:�^���?       ��]�ڕ5@������������������������       �               ;��,��$@�       �                 �u�?��t� �?       ����x&@�       �                 `���?ܗZ�	7�?       i~���@������������������������       �      ȼ       ��/����?������������������������       �               z�5��@������������������������       �               z�5��@������������������������       �               0#0#�?�       �                  �9��?x�d4Fi�??       ���?Y@�       �                 8w�?$�����?       �����8@�       �                 d[�?N��W�?       94���5@�       �                 �ڡ3?�]��0�?       У�Bm�2@�       �                έ���?rR����?       p\����!@�       �                 ��0�?���/��?       U��7�@������������������������       �               �cp>@�       �                   ҏ�?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �               0#0#�?�       �                    �?      �<       /����/#@������������������������       �               ��/���@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               H�4H�4@�       �                 0^�a?R�Q��H�?/       ��nbMS@�       �                 �뜲?g������?       �.�R�3G@�       �                 �Ϻ�?�ң�L��?       ";eQ�<@�       �                  �E�?|��`p��?       �����@������������������������       �               0#0#@������������������������       �      �<       ��/����?�       �                 ��c�?�D��C��?       �c�`�6@������������������������       �               0����/#@�       �                  `���?���6���?       � B��)@�       �                 x��?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#��@�       �                 8Ws�?��d
���?       f�G�N�@������������������������       �               ��/����?�       �                 @B��?;�N9���?       ��{j�@�       �                  ���?��q�R�?       C}Ԥ@�       �                 P�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               0#0# @�       �                  X3�?n��`p��?
       f;3@��1@�       �                 �\��?�;�a
=�?       ��l��@������������������������       �               �cp>@������������������������       �               0#0#�?�       �                   \��?      �<       #0#0&@������������������������       �               0#0# @������������������������       �               vb'vb'"@�       �                 p�B�?�@����?       	}M��=@�       �                  `���?�?�0�!�?       a`�T�4@������������������������       �               0#0#0@�       �                 0���?x�G���?       ��%�|@������������������������       �               0#0# @������������������������       �      �<       ��/����?�       �                    �?hutee�?       Q9��#@������������������������       �               H�4H�4@�       �                 ���?�w��d��?       �0���s@������������������������       �      �<       ��/���@������������������������       �               H�4H�4@�       �                  @���?��1����?0       ��#`T�R@�       �                 @� ?��G�8��?/       v��SR@�       �                  pjS�?B��15�?       ��Qv�-@�       �                 �۶�?���/��?       @z$S��@������������������������       �               ��/����?�       �                 �۲?����?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?�       �                 0��?^����?       �����!@������������������������       �               H�4H�4@�       �                 ����?z��`p��?       �����@������������������������       �               ��/����?������������������������       �      ��       0#0#@�       �                 ����?��I�?"       4j©�,M@�       �                  �Mm�?H�&9���?!       ���ñL@�       �                 �^��?D�r��-�?       ���w�5@�       �                   +Y�?HL�0�h�?       l�e�3@�       �                 ��l�?X�ih�<�?       ��
@������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?������������������������       �      �<       H�4H�4(@�       �                    �?��G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               vb'vb'B@������������������������       �      �<       ��/����?������������������������       �      �<       ��#�� @�t�b��     h�hhK ��h��R�(KK�KK��h �Bx  �k(���e@p�'�x�b@���~�gb@��#��`@��]�ڕU@�A�A.@Np�}^@o��F:lI@H�4H�4@�,����W@�cp>�9@        ��,���A@鰑5@        +�����;@�cp>'@                ��/���@        +�����;@��/���@        *�����;@���-��@        �k(��"@                �k(��2@���-��@        z�5��@���-��@        z�5��@�cp>@                ��/����?        z�5��@��/����?        ;��,��@                ��#���?��/����?                ��/����?        ��#���?                        ��/���@        z�5��(@                        ��/����?        ���>��@/����/#@        z�5��@0����/@        ��#���?��/���@                ��/����?        ��#���?��/����?                ��/����?        ��#���?                ;��,��@��/����?                ��/����?        ;��,��@                ��#���?0����/@        ��#���?                        0����/@        Lp�}N@0����/@        Dy�5A@                �#���9@0����/@        |�5��8@��/����?        z�5��(@��/����?        ;��,��@��/����?        ;��,��@��/����?                ��/����?        ;��,��@                        ��/����?        ���>��@                |�5��(@                ��#���?                [Lg1��&@                ��#���?�cp>@                ��/����?        ��#���?��/����?                ��/����?        ��#���?                z�5��8@��On�8@H�4H�4@;��,��@��|��,@                /����/#@        ;��,��@0����/@        ��#���?��/���@        ��#���?                        ��/���@        ��#��@��/����?                ��/����?        ��#��@                ������3@鰑%@H�4H�4@        �cp>@H�4H�4@        �cp>@0#0#�?        0����/@                ��/����?0#0#�?                0#0#�?        ��/����?                        ��+��+@������3@0����/@        ������3@��/����?        ��#��0@                z�5��@��/����?                ��/����?        z�5��@                        �cp>@        z�5��(@����z�A@vb'vb'"@z�5��(@G�JԮDA@0#0# @z�5��@��/���>@0#0# @z�5��@On��O0@        ��#���?��|��,@                ��|��,@        ��#���?                ;��,��@��/����?        ;��,��@��/����?        ;��,��@                        ��/����?                ��/����?                ��|��,@0#0# @        ��|��,@                        0#0# @z�5��@��/���@        ;��,��@                ��#���?��/���@        ��#���?                        ��/���@                ��/����?�C=�C=@                �C=�C=@        ��/����?        =��,��D@Pn��OP@B�C=ԃ`@�YLg1B@��|��L@^��[�eQ@��b:��:@Nn��O0@��)��)3@z�5��@��/���@��+��+$@        ��/����?        z�5��@��/����?��+��+$@z�5��@��/����?0#0#@        ��/����?0#0#@        ��/����?                        0#0#@z�5��@                                H�4H�4@�,����7@��On�(@vb'vb'"@��#���?�cp>@��+��+@��#���?                        �cp>@��+��+@        �cp>@0#0# @        �cp>@0#0#�?                0#0#�?        �cp>@                ��/����?                ��/����?                        0#0#�?                H�4H�4@[Lg1��6@0����/#@0#0#@        ��/���@        ZLg1��6@�cp>@0#0#@z�5��@��/���@H�4H�4@��#�� @                ��#���?��/���@H�4H�4@��#���?��/���@0#0#�?��#���?        0#0#�?                0#0#�?��#���?                        ��/���@                        0#0# @������3@��/����?0#0#�?������3@��/����?        ;��,��$@                �k(��"@��/����?        z�5��@��/����?                ��/����?        z�5��@                z�5��@                                0#0#�?�k(��"@�)�B�D@l�6k�6I@��#��@���-��*@�C=�C=@��#��@���-��*@0#0#@��#��@���-��*@0#0#�?��#��@��/���@0#0#�?��#��@��/���@                �cp>@        ��#��@��/����?                ��/����?        ��#��@                                0#0#�?        /����/#@                ��/���@                ��/����?                        H�4H�4@                H�4H�4@;��,��@�a#6�;@�
��
�E@;��,��@h
��6@��)��)3@;��,��@On��O0@�C=�C=@        ��/����?0#0#@                0#0#@        ��/����?        ;��,��@��|��,@H�4H�4@        0����/#@        ;��,��@0����/@H�4H�4@��#��@��/����?                ��/����?        ��#��@                ��#���?�cp>@H�4H�4@        ��/����?        ��#���?��/����?H�4H�4@��#���?��/����?0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?��#���?                                0#0# @        �cp>@H�4H�4(@        �cp>@0#0#�?        �cp>@                        0#0#�?                #0#0&@                0#0# @                vb'vb'"@        �cp>@H�4H�48@        ��/����?vb'vb'2@                0#0#0@        ��/����?0#0# @                0#0# @        ��/����?                ��/���@H�4H�4@                H�4H�4@        ��/���@H�4H�4@        ��/���@                        H�4H�4@;��,��@��/���@@�C=�CO@z�5��@��/���@>�C=�CO@z�5��@0����/@�C=�C=@z�5��@�cp>@                ��/����?        z�5��@��/����?        z�5��@                        ��/����?                ��/����?�C=�C=@                H�4H�4@        ��/����?0#0#@        ��/����?                        0#0#@        �cp>@�+��+�K@        ��/����?�+��+�K@        ��/����?��)��)3@        ��/����?vb'vb'2@        ��/����?H�4H�4@                H�4H�4@        ��/����?                        H�4H�4(@        ��/����?0#0#�?                0#0#�?        ��/����?                        vb'vb'B@        ��/����?        ��#�� @                �t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ���JhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKυ�h��BH-         �                 �I�f?�*"��M�?#      ��%	�}@       �                 �^Ҧ?a���w��?�       ���4�xw@       t                 �T�x?"Ik&M��?�       K�����r@       !                  ��?������?�       l��_ik@                        hTl�?��J�s�?       :(']5�E@                        ��;>?��7m�?       �(�+D@                        �ЌT?�Y�t�?       ���bY�@@                           �?�}Cl��?       �(q��;@	                         �!�?�hK)�?       �h��K�2@
                         �fa?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@������������������������       �               ���>��,@                         P�J�?`n����?       ~��Y-"@                        ���R?T����?       P	K��@                          .p�?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@������������������������       �               z�5��@������������������������       �      �<       ��/����?                        @F����/��?       Az$S��@                        0��?Δfm���?       ��Z�N@������������������������       �               ��/����?                         Џ~�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#�� @                        �$I�?      �<       ���-��@������������������������       �               ��/����?������������������������       �               0����/@                         ���?      �<       H�4H�4@������������������������       �               0#0#�?������������������������       �               0#0# @"       ?                 �d�S?�T���?i       _=�y��e@#       .                  �Q�?6�H_�?,       ����L�R@$       '                  @(B�?�y�8��?       47@�=@%       &                  x7?�L����?       Zk���>)@������������������������       �               ��#�� @������������������������       �               鰑%@(       )                  t�޾|M:���?       ����71@������������������������       �               �cp>@*       -                 ���X?\����?	       P	K��,@+       ,                 ��	b?`�s�	�?       f���*@������������������������       �               ��/����?������������������������       �      �<       z�5��(@������������������������       �      ȼ       ��/����?/       >                  lnl?����?       ��y��ZF@0       5                 0��Q?�B���?       �4 �aeE@1       4                    �?���/��?       U��7�@2       3                 �-�?$ k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      �<       ��/���@������������������������       �               z�5��@6       7                 ���	?��i�?       �u�:hA@������������������������       �               ��b:��*@8       ;                    �?�Q0TuJ�?       ȃ�Я[5@9       :                 �4Iw?P�:V��?       �GP�1@������������������������       �        
       ��#��0@������������������������       �      �<       ��/����?<       =                 �)�8?      �<       ��/���@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �      �<       ��/����?@       o                 0�B�?�*.4.�?=       &�)�WY@A       h                 0�2�?L��.�T�?6       es\��V@B       O                    �?B����?.       �R�N�T@C       F                 J�e?�"�d��?       w�I��C@D       E                   ҏ�?
4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @G       L                 ��4�?d!����?       w��^^A@H       I                 ���? �Tu��?       ����>@������������������������       �      ��       �cp>�9@J       K                  �u��?4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @M       N                  �4}?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@P       g                 �jE?h���)�?       �����:E@Q       R                   ��?�I�6��?       �a�ZB@������������������������       �               z�5��@S       Z                 P�p�?X @��?       �\ڞ�@@T       U                 �Sq?�3���r�?       ��7�nN*@������������������������       �               �cp>@V       W                  `���?�FO���?       �ߌ$@������������������������       �      ��       ���>��@X       Y                 �}?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @[       \                  ����?|�b���?       �@cr4@������������������������       �               0����/@]       b                 �=��?z��y�a�?       +��lL/@^       a                 ���?������?       ���'��@_       `                 p���?f%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �               H�4H�4@c       d                 ��?�ۜ�x�?       d��إV#@������������������������       �               ��/���@e       f                 �[�Z?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               �cp>@i       l                 /0�?8�j���?       ���z"@j       k                  ��ľ      �<       ���>��@������������������������       �               ;��,��@������������������������       �               ��#�� @m       n                 ����?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?p       s                 �K��?p@����?       ���a�#@q       r                  �"�?d*�'=P�?        �2"@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      ȼ       ��/����?u       ~                      ���^�?-       bʂM,�S@v       {                  ��?�CPͳ�?       �I6��B@w       x                    �?��+�*�?       yȚ�
A@������������������������       �        
       ������3@y       z                     �?H�=�Sο?       ����,@������������������������       �               ��/����?������������������������       �      ��
       ��b:��*@|       }                  0B�?���`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @       �                  ���?$���~D�?       �ܻd؂D@�       �                 @�_�?d�WT�V�?	       C$_]3@�       �                 @��?�C=+��?       b��T|0@������������������������       �      ��       ���>��,@�       �                 sT�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 (�S?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?�       �                    �?��_~"��?       �bj��5@�       �                 ��8�?nQ��?
       �s�=�1@������������������������       �      ��       ��On�(@�       �                 �q�?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?�       �                 ��K�? �J���?       ��*]Y@������������������������       �               0#0# @������������������������       �               ��#�� @�       �                 �%��?��!a�w�?5       r����S@�       �                 P�8�?N*�<��?       �"3���E@�       �                  �u��?��r�S�?       �f��%/@�       �                 � ��?e��}�?
       ��Se+@�       �                  ���?$ k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      ��       ��/���@�       �                 ���?      �<       E�JԮD!@������������������������       �               ��/����?������������������������       �               ��/���@������������������������       �               0#0# @�       �                  �d%�? 2�x^�?       ���,$�;@�       �                 0�ݮ?��G�%�?       \��rs2@������������������������       �               H�4H�4@�       �                 pHF�?�Tu��?       ����.@�       �                 �[��?$ k�Lj�?       �q��l}@������������������������       �      ��       �cp>@�       �                �ܷB�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 ���@?      �<       鰑%@������������������������       �               /����/#@������������������������       �               ��/����?������������������������       �               vb'vb'"@�       �                ����}?�����?       ���7~�A@�       �                 �Y|�?pa��6��?       ���$@4@�       �                 ����?�|2N��?       �3K}@������������������������       �               0#0#�?�       �                 �QT�?�zœ���?       IG���t@������������������������       �               z�5��@������������������������       �               0#0#�?������������������������       �        
       �A�A.@�       �                 �N��?=!eM-f�?	       �L+��-@������������������������       �               H�4H�4@�       �                 0ֺ�?�C>�?       �1�m�!@������������������������       �               �cp>@�       �                 ����?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?�       �                    �?|����?@       Xy��+ X@�       �                 ��?YG篓�?        ��:I@������������������������       �               ��#���?������������������������       �               [��Y��H@�       �                 @F�`��8���?        �cp>G@������������������������       �               ��/����?�       �                 ��e�?�q��/��?       h
��F@�       �                 ��N�?�:�^���?       ��]�ڕE@�       �                 )��?��i���?       ����A@�       �                 ��;�?�-�bƲ?       >�7*9@������������������������       �               H�4H�48@������������������������       �      �<       ��/����?�       �                 �?���`p��?       f;3@��!@�       �                  �Ԧ�?�@G���?       hu��@�       �                 ���?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 �p�?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��+��+@������������������������       �               vb'vb'"@������������������������       �      �<       ��/����?�t�bh�hhK ��h��R�(KK�KK��h �Bh  ?��,��d@D:l��d@}��z�Gb@-�����d@.����/c@�[��[�L@������c@2��18^@��)��)3@�5��P�Y@k��F:lY@�A�A.@��b:��:@���-��*@H�4H�4@��b:��:@���-��*@        ��b:��:@���-��@        �,����7@��/���@        ��,���1@��/����?        z�5��@��/����?                ��/����?        z�5��@                ���>��,@                z�5��@�cp>@        z�5��@��/����?        z�5��@��/����?                ��/����?        z�5��@                z�5��@                        ��/����?        z�5��@�cp>@        ��#���?�cp>@                ��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#�� @                        ���-��@                ��/����?                0����/@                        H�4H�4@                0#0#�?                0#0# @B����R@h
��V@H�4H�4(@5��tSH@�cp>�9@        ���>��,@��/���.@        ��#�� @鰑%@        ��#�� @                        鰑%@        z�5��(@0����/@                �cp>@        z�5��(@��/����?        z�5��(@��/����?                ��/����?        z�5��(@                        ��/����?        Ey�5A@鰑%@        Ey�5A@D�JԮD!@        ��#��@��/���@        ��#���?��/���@        ��#���?                        ��/���@        z�5��@                Jp�}>@0����/@        ��b:��*@                ��#��0@0����/@        ��#��0@��/����?        ��#��0@                        ��/����?                ��/���@                ��/����?                ��/����?                ��/����?        ��b:��:@3����-O@H�4H�4(@��b:��:@=��18N@0#0#@�k(��2@�_��e�M@0#0#@��#��@F�JԮDA@0#0#�?��#�� @�cp>@                �cp>@        ��#�� @                ��#�� @�]�ڕ�?@0#0#�?��#�� @��|��<@                �cp>�9@        ��#�� @�cp>@                �cp>@        ��#�� @                        �cp>@0#0#�?                0#0#�?        �cp>@        ���>��,@��On�8@H�4H�4@���>��,@0����/3@H�4H�4@z�5��@                [Lg1��&@0����/3@H�4H�4@�k(��"@��/���@                �cp>@        �k(��"@��/����?        ���>��@                ��#�� @��/����?                ��/����?        ��#�� @                ��#�� @��/���.@H�4H�4@        0����/@        ��#�� @鰑%@H�4H�4@��#���?��/����?H�4H�4@��#���?��/����?                ��/����?        ��#���?                                H�4H�4@��#���?D�JԮD!@                ��/���@        ��#���?��/����?                ��/����?        ��#���?                        �cp>@        ��#�� @��/����?        ���>��@                ;��,��@                ��#�� @                ��#���?��/����?                ��/����?        ��#���?                        ��/����?0#0# @        ��/����?0#0# @        ��/����?                        0#0# @        ��/����?        �>��nK@/����/3@0#0#@��#��@@��/����?0#0# @��#��@@��/����?        ������3@                ��b:��*@��/����?                ��/����?        ��b:��*@                        ��/����?0#0# @        ��/����?                        0#0# @�k(���5@E�JԮD1@0#0# @�P^Cy/@��/���@        �P^Cy/@��/����?        ���>��,@                ��#���?��/����?        ��#���?                        ��/����?                �cp>@                ��/����?                ��/����?        z�5��@���-��*@0#0# @��#��@���-��*@                ��On�(@        ��#��@��/����?        ��#��@                        ��/����?        ��#�� @        0#0# @                0#0# @��#�� @                ���>��@Pn��O@@��)��)C@��#�� @���-��:@�C=�C=,@��#���?��On�(@0#0# @��#���?��On�(@        ��#���?��/���@        ��#���?                        ��/���@                E�JԮD!@                ��/����?                ��/���@                        0#0# @��#���?��|��,@H�4H�4(@��#���?��|��,@H�4H�4@                H�4H�4@��#���?��|��,@        ��#���?��/���@                �cp>@        ��#���?��/����?                ��/����?        ��#���?                        鰑%@                /����/#@                ��/����?                        vb'vb'"@;��,��@�cp>@H�4H�48@z�5��@        S2%S2%1@z�5��@        0#0# @                0#0#�?z�5��@        0#0#�?z�5��@                                0#0#�?                �A�A.@��#�� @�cp>@�C=�C=@                H�4H�4@��#�� @�cp>@0#0#�?        �cp>@        ��#�� @        0#0#�?��#�� @                                0#0#�?��#���?���-��@#0#0V@��#���?        \��Y��H@��#���?                                [��Y��H@        ���-��@������C@        ��/����?                0����/@������C@        ��/���@������C@        ��/���@�A�A>@        ��/����?H�4H�48@                H�4H�48@        ��/����?                �cp>@H�4H�4@        �cp>@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?                ��/����?                ��/����?                        ��+��+@                vb'vb'"@        ��/����?        �t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�
HyhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKㅔh��B�1         �                 0�0�?֗�O�?+       0۽�v}@       �                 ����?*w��J�?�       �}�3��s@       ~                 в��?1j��rs�?�       �5��"q@                        ����?�*��Q��?�       h�3"Y�o@                        �UH{?`$�*��?       N{���2@                        0��?�4��v�?       �Y-"�'@������������������������       �               ��/���@                         ��^�?>9�)\e�?       _���b @	       
                 `��$?
4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @������������������������       �               z�5��@                        b?X�ih�<�?       ��
@                        �G��?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �      ��       H�4H�4@       A                 �o?�p>�])�?�       �b1�Im@       (                  _z_?�iφ�z�??       �n�>%�Z@       %                 @Ws�?^dؗ��?       4d��8@       "                 `%�7?* k�Lj�?       �q��l}3@                        P���>��|��?
       ���ĺw+@������������������������       �               �cp>@                        �$?Z?���3�?	       ���(+�%@                        p��I?dQ��?       �s�=�!@������������������������       �               ��#���?                        ��^^?l�r{��?       e�6� @������������������������       �               �cp>@                         9U?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?        !                  �~��?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?#       $                   ���?      �<       �cp>@������������������������       �               �cp>@������������������������       �               �cp>@&       '                    �?ܗZ�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@)       4                 �|y?vM��vn�?/       ���eA�T@*       3                 ��8�?X#W�+�?       �W�EaD@+       ,                  Pmj�?X
TI
u�?       �إV�C@������������������������       �               ��/����?-       0                  qUi?��p?��?       P�^��B@.       /                 ��%f?�FO���?       �ߌ$@������������������������       �      ��       �k(��"@������������������������       �      ȼ       ��/����?1       2                 @F�      �<       ��b:��:@������������������������       �               :��,��4@������������������������       �               z�5��@������������������������       �      �<       ��/����?5       >                 @*tC?�)z� ��?       a��!E@6       =                 `�ג?�M:���?       ����7A@7       8                 ��$?x�n3��?       ƛ2��4@������������������������       �               �k(��"@9       :                  �.þt@ȱ��?       nm���S'@������������������������       �      ��       D�JԮD!@;       <                 0?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �        	       ��b:��*@?       @                  9�>      �<       ��/���@������������������������       �               �cp>@������������������������       �               0����/@B       E                  h��?<��k�f�?M        W֏��_@C       D                 �/��?b,���O�?       ���/>@������������������������       �               ��#���?������������������������       �               H�4H�4@F       i                 ��\�?������?J       �����^@G       ^                 `��g?�l?�07�?1       �u��-S@H       [                  T?2��n��?       ]����H@I       Z                 @j��?䶎�h�?       ���9�E@J       M                    �?h~p �?       ���!�DE@K       L                 `U�?      �<       �e�_��7@������������������������       �               �cp>'@������������������������       �               ��On�(@N       O                 芋�?F�tg��?       c�㡍2@������������������������       �               ��/���@P       Q                 �k?�!�GU�?       m�����%@������������������������       �               ��#�� @R       U                 PU1�?�`���6�?       /u��֝!@S       T                 ��z�?      �<       ��/���@������������������������       �               ��/����?������������������������       �               �cp>@V       W                 �p�?��`i��?       �؛.�@������������������������       �               0#0# @X       Y                 ����?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      �<       ��#���?\       ]                 p'v�?ln����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#��@_       f                  Q��?v���E`�?       s��u;@`       c                 0�{?T�'e��?       �F�ҽn0@a       b                 `|��?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @d       e                 TVT?T�s�	�?       e���*@������������������������       �               z�5��(@������������������������       �      ȼ       ��/����?g       h                 �s$�?��XnP��?       ѭS`oM%@������������������������       �               E�JԮD!@������������������������       �               0#0# @j       w                 ��{�?��*P���?       �	�kjG@k       r                 0�2�?,�D��?       �>Dq6/=@l       m                 t��t? �w�]��?       !5��o�/@������������������������       �               ��/���@n       q                 ��.�?��<��?       t=�x�(@o       p                 p�T�?��6L�n�?       �E#��h @������������������������       �      �<       ���>��@������������������������       �      ȼ       ��/����?������������������������       �      м       ��/���@s       v                 ����?�(߫$��?       2H����*@t       u                    �?      �<       [Lg1��&@������������������������       �               ���>��@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?x       y                 @U�?��/ʪ��?       H�Ų��1@������������������������       �               z�5��@z       {                 ��?|���A�?	       /gX\-@������������������������       �               ��/���@|       }                 ����?��|��?       ���ĺw@������������������������       �               0����/@������������������������       �               ��#�� @       �                 ��]�?Bv��l��?       ���Q��4@�       �                 ����?ǳ�F�M�?       S��ڭQ(@������������������������       �               H�4H�4@�       �                 �a��?"�wO��?       ����D"@������������������������       �               0#0# @�       �                 �ߦx?|��j�?       �e��w@�       �                    �?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �               0#0# @�       �                  y��?�`���6�?       .u��֝!@������������������������       �               0#0# @�       �                 �ڽ?�`@s'��?       Ei_y,*@������������������������       �               ��#���?������������������������       �               �cp>@�       �                  X?�Y}��K�?       `��D@�       �                �S�|?~�[����?       ^~.1<@�       �                 0��?��Vj��?       s�{R�:@�       �                  @���?�T�V���?       �a���!2@�       �                   .p�?�6��b�?       %�|�1@������������������������       �               ��/����?������������������������       �      ��
       0#0#0@������������������������       �      �<       ��#���?�       �                 �m��?����|e�?       �z �B�@������������������������       �               H�4H�4@�       �                 �/�?lutee�?       Q9��@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                 �s�?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?�       �                 �l��?      �<	       H�4H�4(@������������������������       �               0#0#�?������������������������       �               #0#0&@�       �                 �Y8�?[]߆B�?h       _d�y�c@�       �                 �b'�?�x�PX�?)       �:�,0Q@�       �                  ���?��3v���?       l�--��8@�       �                 �zm�?|�و��?       bR4��/@�       �                 p�v�?�AP�9��?       i��6��@������������������������       �               0#0#@�       �                  ���?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 �u�b?�`���6�?       /u��֝!@�       �                 8*��?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?�       �                 P���?<�a
=�?       ��l��@������������������������       �               0����/@�       �                 �yo�?z�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               vb'vb'"@�       �                 �Y�?�o����?       ޞ�3��E@�       �                 ���l?�:�D���?       b�V�RlB@�       �                  �^��?X�s�	�?       f���:@������������������������       �               ��/����?�       �                 ��ߞ?���OT�?       p�>%,�9@������������������������       �               ��/����?������������������������       �               z�5��8@�       �                 `&�?      �<       ��+��+$@������������������������       �               0#0# @������������������������       �               0#0# @������������������������       �      м       �C=�C=@�       �                 ��u�?h��ߗ��??       �D�V@�       �                 p&�?�:g�Q�?       ��ʭ�0@������������������������       �               0#0# @�       �                 �6�?���p�?       f-��VS-@�       �                 �d��?p .A��?       �wPq�@������������������������       �               �cp>@�       �                 �؉�?�o���?       o�9�F@������������������������       �               0#0#@������������������������       �               ��#���?������������������������       �      ��       ���-��@�       �                 �'٪?6�T_��?1       �D�XB�Q@�       �                  �E�?�P�`B�?	       �F�N@�0@�       �                 ��ǻ?�֪u�_�?       ��?�8'@�       �                 �$I�?|�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      ��       ��/���@������������������������       �               ��+��+@�       �                 ����?��g����?(       �f��K@�       �                 �qҍ?�u�����?'       6�6�K@�       �                  ~�?�N�����?       �j4�M�;@�       �                 @�-�?|�G���?       ��%�|/@�       �                 ����?�v�;B��?       ՟���	 @������������������������       �               ��/����?������������������������       �               �C=�C=@�       �                 �ʎ�?xLU���?       h�ҹ^�@������������������������       �               ���-��@������������������������       �               0#0#�?�       �                  <�?T������?	       "�B(@������������������������       �               �C=�C=@�       �                  ��?�o���?       o�9�F@������������������������       �               ��#���?������������������������       �               0#0#@�       �                  0@�?      �<       ��8��8:@������������������������       �               0#0#�?������������������������       �               k�6k�69@������������������������       �      �<       ��/����?�t�bh�hhK ��h��R�(KK�KK��h �BH  y�YLGc@]�ڕ��d@�����b@'�}��_@n>�c0`@�s?�s?M@	�#�O_@(����-_@H�4H�48@Np�}^@�����]@�A�A.@;��,��@��/���@H�4H�4@;��,��@���-��@                ��/���@        ;��,��@�cp>@        ��#�� @�cp>@                �cp>@        ��#�� @                z�5��@                        ��/����?H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@                H�4H�4@��P^C�\@M!Д[@vb'vb'"@Fy�5Q@2����/C@        ���>��@E�JԮD1@        ��#��@��/���.@        ��#��@/����/#@                �cp>@        ��#��@���-��@        ��#�� @���-��@        ��#���?                ��#���?���-��@                �cp>@        ��#���?��/����?                ��/����?        ��#���?                ��#�� @                ��#���?                ��#���?                        �cp>@                �cp>@                �cp>@        z�5��@��/����?                ��/����?        z�5��@                ��>���N@鰑5@        �YLg1B@��/���@        �YLg1B@��/����?                ��/����?        �YLg1B@��/����?        �k(��"@��/����?        �k(��"@                        ��/����?        ��b:��:@                :��,��4@                z�5��@                        ��/����?        z�5��8@D�JԮD1@        {�5��8@/����/#@        [Lg1��&@0����/#@        �k(��"@                ��#�� @0����/#@                D�JԮD!@        ��#�� @��/����?        ��#�� @                        ��/����?        ��b:��*@                        ��/���@                �cp>@                0����/@        ����JG@����Q@vb'vb'"@��#���?        H�4H�4@��#���?                                H�4H�4@]Lg1��F@����Q@H�4H�4@�k(���5@y%jW�vH@H�4H�4@��#�� @������C@0#0# @��#��@�+Q��B@0#0# @z�5��@�+Q��B@0#0# @        �e�_��7@                �cp>'@                ��On�(@        z�5��@���-��*@0#0# @        ��/���@        z�5��@�cp>@0#0# @��#�� @                ��#���?�cp>@0#0# @        ��/���@                ��/����?                �cp>@        ��#���?��/����?0#0# @                0#0# @��#���?��/����?        ��#���?                        ��/����?        ��#���?                ��#��@��/����?                ��/����?        ��#��@                ��b:��*@0����/#@0#0#@��b:��*@��/����?0#0# @��#���?        0#0# @��#���?                                0#0# @z�5��(@��/����?        z�5��(@                        ��/����?                E�JԮD!@0#0# @        E�JԮD!@                        0#0# @�,����7@�cp>7@        �k(��2@鰑%@        ���>��@D�JԮD!@                ��/���@        ���>��@0����/@        ���>��@��/����?        ���>��@                        ��/����?                ��/���@        ZLg1��&@��/����?        [Lg1��&@                ���>��@                ��#��@                        ��/����?        ;��,��@��On�(@        z�5��@                ��#�� @��On�(@                ��/���@        ��#�� @0����/@                0����/@        ��#�� @                ;��,��@���-��@vb'vb'"@��#��@��/����?�C=�C=@                H�4H�4@��#��@��/����?0#0#@                0#0# @��#��@��/����?0#0# @��#��@��/����?                ��/����?        ��#��@                                0#0# @��#���?�cp>@0#0# @                0#0# @��#���?�cp>@        ��#���?                        �cp>@        ��#���?0����/@T2%S2%A@��#���?0����/@#0#06@��#���?�cp>@#0#06@��#���?��/����?0#0#0@        ��/����?0#0#0@        ��/����?                        0#0#0@��#���?                        ��/����?H�4H�4@                H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@        ��/����?                ��/����?                ��/����?                        H�4H�4(@                0#0#�?                #0#0&@*�����;@�+Q��B@ �q��V@�#���9@0����/#@B�A�@@��#���?��/���@0#0#0@��#���?��/���@�C=�C=@        ��/����?��+��+@                0#0#@        ��/����?0#0#�?                0#0#�?        ��/����?        ��#���?�cp>@0#0# @��#���?        0#0#�?��#���?                                0#0#�?        �cp>@0#0#�?        0����/@                ��/����?0#0#�?                0#0#�?        ��/����?                        vb'vb'"@z�5��8@��/����?S2%S2%1@{�5��8@��/����?��+��+$@z�5��8@��/����?                ��/����?        z�5��8@��/����?                ��/����?        z�5��8@                                ��+��+$@                0#0# @                0#0# @                �C=�C=@��#�� @�a#6�;@�s?�s?M@��#���?0����/#@H�4H�4@                0#0# @��#���?0����/#@0#0#@��#���?�cp>@0#0#@        �cp>@        ��#���?        0#0#@                0#0#@��#���?                        ���-��@        ��#���?;l��F:2@��8��8J@        /����/#@�C=�C=@        0����/#@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @        ��/���@                        ��+��+@��#���?D�JԮD!@;�;�F@��#���?��/���@;�;�F@��#���?��/���@��)��)3@        ��/���@0#0# @        ��/����?�C=�C=@        ��/����?                        �C=�C=@        ���-��@0#0#�?        ���-��@                        0#0#�?��#���?        #0#0&@                �C=�C=@��#���?        0#0#@��#���?                                0#0#@                ��8��8:@                0#0#�?                k�6k�69@        ��/����?        �t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ���]hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK߅�h��B�0         �                 �8��?�'�ѧK�?0      ���P>�}@       w                   ��?���J�?�       �m��+�s@       d                 �&�?��쑎�?�       �҇M+o@       9                 `=&�?w)�8�^�?�       Ȳ{H~j@       0                 ��??
e���?Y       8����a@       -                  ���? M����?C       +#߫�"\@                        �C
T?�RQHB�?>       �\S'y�Y@                        ,*����\#�C�?        2`R;J@	                        09h? Z��K�?       ��K�M�:@
                        �&�?���/��?       ���U�5@                        N��S?��߭Q��?
       �QVl�0@                        � Q	?4=�%�?        t=�x�-@                        �-�?�PJo�x�?       T|qt�&@������������������������       �               �cp>@                         �.�?����?       ��X�)B @������������������������       �               ��/����?������������������������       �      �<       z�5��@������������������������       �      м       ��/���@������������������������       �               ��/����?������������������������       �      �<       ;��,��@                        �N-?     ��<       0����/@������������������������       �               ��/����?������������������������       �               ��/���@                        ��X?���P��?       �*Y�ȹ9@������������������������       �               ��/����?������������������������       �      �<       �,����7@       &                 ����?<��s��?       �XT>�!I@       !                   s��?��y6t�?       E�RN��C@                        ��py?���m�?       .���<@������������������������       �               <��,��4@                         `�?��6L�n�?       �E#��h @������������������������       �               ��/����?������������������������       �      �<       ���>��@"       #                  ��d�?�d�$���?       �T�f$@������������������������       �               ��/����?$       %                    �?      �<       ��#�� @������������������������       �               ;��,��@������������������������       �               z�5��@'       ,                  �j?���Ѯ�?       ��GQ&@(       +                   \��?�d�$���?       �T�f$@)       *                ���[�?      �<       ��#�� @������������������������       �               ��#��@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �      м       ��/����?.       /                 {X?������?       �4^$4�#@������������������������       �               z�5��@������������������������       �               ���-��@1       8                  gm?ar[+Z�?       
i!�Y<@2       5                  ����?LG�:">�?       �K��G:@3       4                 H���?@H�,.̷?       �J�$r.5@������������������������       �               &jW�v%4@������������������������       �      �<       ��#���?6       7                 h�B?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �      �<       ��#�� @:       Q                 ����?��>s��?)       �),��Q@;       <                 ����?`sm+�?       W�|���A@������������������������       �               �C=�C=@=       >                 �`?���p���?       ���� r<@������������������������       �               0#0# @?       J                 �$܀?$��	�C�?       q_��m:@@       A                 �-�~?�p���K�?       D2(ߪ{0@������������������������       �               D�JԮD!@B       I                XI
|�?���`�?       ��
�Me@C       H                  ����?��n��?       �-H�\@D       G                 ��=�?��q�R�?       C}Ԥ@E       F                  pjS�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �      ��       ��/���@������������������������       �               0#0#�?K       P                 �~N?��
+���?       \Zz�+�#@L       M                    �?�djH�E�?       ^�\m�n@������������������������       �               ��#��@N       O                 p���?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       ��/���@R       S                 �it?rsxI�?       ���r�A@������������������������       �               �cp>@T       c                 �p�?��M��?       W��%U@@U       X                  ��?䪃�h��?       ��(�?@V       W                 ��;�?& k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      �<       ��/���@Y       Z                 ����?�F�o��?       '��:@������������������������       �               �P^Cy/@[       \                 �2*�?�w�ٕ��?       sǩ���&@������������������������       �               0#0# @]       `                  �5�?X�j���?       ���z"@^       _                 0�qw?����?       ��X�)B@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?a       b                 ��N�?      �<       ;��,��@������������������������       �               ��#���?������������������������       �               ��#��@������������������������       �               0#0#�?e       r                 ���?� ���+�?       �+TG�B@f       g                  .z�?��_.���?       ��C��>@������������������������       �               0#0# @h       i                 �o��?nw��?       c�?�-<@������������������������       �               h
��6@j       k                 x��?��q�R�?       C}Ԥ@������������������������       �               0#0# @l       q                  ZeK?���/��?       V��7�@m       n                  mI�?`n����?       � ��w<@������������������������       �               ��#���?o       p                 ��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      �<       ��/����?s       t                 X�)�?0y��]0�?       ���y"@������������������������       �               0#0#@u       v                 (o�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?x       �                 д��?d�P�a��?%       ��oW*P@y       z                 0��?���A���?       ��\�F2@������������������������       �               ��/����?{       �                 �5�?v�w�o�?       �c/�P1@|                        @�0?�~�Hs=�?       ��?Z[0@}       ~                 ��7�?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?�       �                 �A�?��ڰ�x�?
       �K�f�(@������������������������       �        	       <��,��$@������������������������       �               0#0# @������������������������       �      �<       ��/����?�       �                 P���?�����?       ���i1G@�       �                  �<F?�Y�R���?       v��\�A@�       �                 0��?���1p8�?       |곯�+@�       �                 �-�?f%@�"�?       ��[�@������������������������       �      �<       ��/���@������������������������       �               ��#�� @������������������������       �               0#0# @������������������������       �      ��       ��-��-5@�       �                 �fQ?d�wy��?       �f0�v&@�       �                  `%+�?��6L�n�?       �E#��h @������������������������       �               ��#��@�       �                 ���?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@������������������������       �               H�4H�4@�       �                 p- �?�p���m�?o       �G�%�c@�       �                  `��?�����?       ޕ:��|>@�       �                 ��v�?��E9p5�?       s4agv;@�       �                 ����?Dm����?       ��?��7@�       �                    �?�a����?
       
AC6&@������������������������       �               ;��,��@�       �                 `Ձ�?vT �+��?       ��>Y��@�       �                ��r�?Ȕfm���?       ��Z�N@������������������������       �               ��#���?�       �                 H8��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               0#0# @�       �                 �3��?x�+%�"�?       ��kw��(@������������������������       �      ��       [Lg1��&@������������������������       �               0#0#�?�       �                 ��(�?H��NV=�?       �t�ܲ@������������������������       �               ��/����?�       �                 �Dr�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               H�4H�4@�       �                 �cp�?�c��@�?Y       ����.`@�       �                 Ў m?!&k���?=       �ё,��V@�       �                 ��{�?�V���?       ���F@�       �                 �D��?����|e�?       �z �B�@������������������������       �               ��+��+@�       �                 ��8�?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?�       �                 �I�?�8vfd�?       h��\��B@�       �                 ���D?ڭ�8&S�?       �x��T&?@�       �                 �b'�?��t?��?       "���5�3@������������������������       �               0#0# @�       �                 �!�?���;�1�?       �$�S՞1@�       �                 06Υ?��c`�?       %��t5)@������������������������       �               ��#���?������������������������       �               �cp>'@�       �                  �?�nɵ��?       Cad�J@�       �                 �^��?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �      ��       z�5��@�       �                 �T�?      �<	       �cp>'@������������������������       �               ��/����?������������������������       �               鰑%@�       �                    �?ln����?       � ��w<@�       �                 ��޴?`%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               z�5��@�       �                 �'m�?�o�k��?       4���G@�       �                    �?�8M�ҿ?       .2�&�E@������������������������       �               ��+��+4@�       �                  `�J�? ��q��?       �?8��7@������������������������       �               H�4H�4(@�       �                 XR��?���};��?	       ��;̑�%@�       �                  `%+�?~�G���?       '5L�`�@������������������������       �               �cp>@������������������������       �               H�4H�4@������������������������       �               ��+��+@�       �                p���? �� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 pg_�?�?�	,�?       ?0�1bC@�       �                 ��X�?�=�
��?       o��V��6@�       �                  �~��?H,�#6?�?       ���*4@�       �                 �=��?Hy��]0�?       ���y"@������������������������       �               ��/����?������������������������       �               ��+��+@������������������������       �      ��       �C=�C=,@�       �                 �?�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?�       �                 ��F�?      �<       �A�A.@������������������������       �               0#0# @������������������������       �               ��8��8*@�t�bh�hhK ��h��R�(KK�KK��h �B�  ��P^CYe@q�'�x�b@�����b@�}��a@M!Д[@�s?�s?M@��>���^@l��F:lY@H�4H�48@Np�}^@3����/S@�A�A.@:��P^�V@q��F:lI@        >��,��T@�_��e�=@        �b:���S@�cp>7@        ��,���A@E�JԮD1@        ZLg1��&@��/���.@        ZLg1��&@鰑%@        z�5��@鰑%@        z�5��@E�JԮD!@        z�5��@0����/@                �cp>@        z�5��@��/����?                ��/����?        z�5��@                        ��/���@                ��/����?        ;��,��@                        0����/@                ��/����?                ��/���@        �,����7@��/����?                ��/����?        �,����7@                �GpAF@�cp>@        �YLg1B@�cp>@        )�����;@��/����?        <��,��4@                ���>��@��/����?                ��/����?        ���>��@                ��#�� @��/����?                ��/����?        ��#�� @                ;��,��@                z�5��@                ��#�� @�cp>@        ��#�� @��/����?        ��#�� @                ��#��@                ��#��@                        ��/����?                ��/����?        z�5��@���-��@        z�5��@                        ���-��@        ���>��@鰑5@        ;��,��@鰑5@        ��#���?&jW�v%4@                &jW�v%4@        ��#���?                ��#��@��/����?                ��/����?        ��#��@                ��#�� @                Jp�}>@�cp>�9@�A�A.@;��,��@:l��F:2@H�4H�4(@                �C=�C=@;��,��@;l��F:2@��+��+@                0#0# @;��,��@9l��F:2@H�4H�4@��#���?���-��*@0#0# @        D�JԮD!@        ��#���?0����/@0#0# @��#���?0����/@0#0#�?��#���?��/����?0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?��#���?                        ��/���@                        0#0#�?��#��@0����/@0#0#�?��#��@��/����?0#0#�?��#��@                        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/���@        {�5��8@��/���@H�4H�4@        �cp>@        {�5��8@0����/@H�4H�4@{�5��8@0����/@0#0# @��#���?��/���@        ��#���?                        ��/���@        �,����7@��/����?0#0# @�P^Cy/@                ��#�� @��/����?0#0# @                0#0# @��#�� @��/����?        z�5��@��/����?        z�5��@                        ��/����?        ;��,��@                ��#���?                ��#��@                                0#0#�?��#�� @��On�8@vb'vb'"@��#�� @�e�_��7@0#0#@                0#0# @��#�� @�e�_��7@0#0# @        h
��6@        ��#�� @��/����?0#0# @                0#0# @��#�� @��/����?        ��#�� @��/����?        ��#���?                ��#���?��/����?        ��#���?                        ��/����?                ��/����?                ��/����?��+��+@                0#0#@        ��/����?0#0#�?        ��/����?                        0#0#�?�k(���5@D�JԮD!@S2%S2%A@|�5��(@��/���@0#0# @        ��/����?        |�5��(@�cp>@0#0# @|�5��(@��/����?0#0# @��#�� @��/����?        ��#�� @                        ��/����?        <��,��$@        0#0# @<��,��$@                                0#0# @        ��/����?        �k(��"@0����/@0#0#@@��#�� @��/���@�s?�s?=@��#�� @��/���@0#0# @��#�� @��/���@                ��/���@        ��#�� @                                0#0# @                ��-��-5@���>��@��/����?H�4H�4@���>��@��/����?        ��#��@                z�5��@��/����?                ��/����?        z�5��@                                H�4H�4@��b:��:@�)�B�D@"�q��V@�k(��2@0����/@�C=�C=@�k(��2@0����/@0#0#@��,���1@�cp>@H�4H�4@z�5��@�cp>@0#0# @;��,��@                ��#���?�cp>@0#0# @��#���?�cp>@        ��#���?                        �cp>@                ��/����?                ��/����?                        0#0# @[Lg1��&@        0#0#�?[Lg1��&@                                0#0#�?��#���?��/����?0#0#�?        ��/����?        ��#���?        0#0#�?��#���?                                0#0#�?                H�4H�4@��#�� @;l��F:B@��-��-U@��#�� @On��O@@n�6k�6I@��#�� @�a#6�;@vb'vb'"@        ��/����?H�4H�4@                ��+��+@        ��/����?0#0#�?        ��/����?                        0#0#�?��#�� @�cp>�9@H�4H�4@��#��@�e�_��7@H�4H�4@��#��@��On�(@H�4H�4@                0#0# @��#��@��On�(@0#0#�?��#���?�cp>'@        ��#���?                        �cp>'@        z�5��@��/����?0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?        z�5��@                        �cp>'@                ��/����?                鰑%@        ��#��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        z�5��@                        0����/@�ڬ�ڬD@        �cp>@��+��+D@                ��+��+4@        �cp>@��+��+4@                H�4H�4(@        �cp>@0#0# @        �cp>@H�4H�4@        �cp>@                        H�4H�4@                ��+��+@        ��/����?0#0#�?                0#0#�?        ��/����?                ��/���@S2%S2%A@        ��/���@��)��)3@        ��/����?��)��)3@        ��/����?��+��+@        ��/����?                        ��+��+@                �C=�C=,@        �cp>@                ��/����?                ��/����?                        �A�A.@                0#0# @                ��8��8*@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�;hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK���h��B6         �                 �=��?�i�TpQ�?-      Me=�w}@       �                  �=�?f�����?�       P(!EDw@       �                 �I�f?�	m�{�?�       ����p@       A                 0%�z?Ӂ��ӏ�?�       ��'Х*n@       6                 �:W>?X�M5^�?H       [�׭-?[@                        �U����,A���??       ++�aW@                        ��V?��`;�?       �N��?C@                         `<��?nQ��?       �s�=�!@	       
                 h�[�>�`@s'��?       Fi_y,*@������������������������       �               ��#���?                        �?9?      �<       �cp>@������������������������       �               ��/����?������������������������       �               0����/@                        HԱ?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?                        ��V?��{�b��?       zc�)ai=@                          �P�?�4��v�?       �Y-"�'@                        G+�`?� �_rK�?       J�@��"@                         �g<�?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �      ��       ��#��@                         �"�?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �      ȼ       �cp>@                         �G?�?x�:V��?       �GP�1@������������������������       �               ��/����?������������������������       �               ��#��0@       '                 ���#?Ɣr��%�?$       �z��K@       $                 ���p?h7uV��?       m}�'�:@        #                  �6�?�����?       �O��@!       "                 �Q�?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               z�5��@%       &                    �?      �<       <��,��4@������������������������       �        	       ���>��,@������������������������       �               z�5��@(       3                  P�"�?��h!��?       [�v%jW;@)       .                    �?^�T��?       ��R�)@*       -                  �я�?h�r{��?       e�6� @+       ,                 P�2?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               ��/���@/       2                 `%�7?�d�$���?       �T�f@0       1                 �R�*?      �<       ��#��@������������������������       �               ��#�� @������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?4       5                    �?      �<
       ���>��,@������������������������       �        	       ��b:��*@������������������������       �               ��#���?7       <                 ����?�(�����?	       ��0��0@8       ;                 �<�?�F���?       :�.�-'@9       :                 Y]?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �               E�JԮD!@=       >                 `�??�Z�	7�?       j~���@������������������������       �               ��#�� @?       @                 h�� ?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?B       w                  `���?�x����?V       ��;��`@C       p                 ГӢ?Σ^�hl�?A       /�g�X@D       U                 �}�Y?�},p�?8       �Ք%�U@E       T                 ��_�?����w�?       ���Ã@?@F       M                 �1�?$#�-�?       ��$=�%<@G       L                 �Н�?�^�#΀�?       O�{��A5@H       I                 �-�?��٤ݸ?       ��<5�84@������������������������       �               �cp>'@J       K                  h?)���?       y��uk!@������������������������       �               ��#���?������������������������       �               ��/���@������������������������       �      �<       ��#���?N       O                 �%s?l��w��?       ���@������������������������       �               ��#���?P       S                  �Q�?�� ��?       qp� k@Q       R                 M_?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               �cp>@������������������������       �      ȼ       z�5��@V       o                 `��?H��I��?$       kF�G	�K@W       j                 �?�4�8��?#       ��`�7J@X       g                 �,�?�Ug���?       ����@@Y       `                 Pz�?`�T��?       ��R�9@Z       _                 TVT?��?       ��l}�'*@[       \                 �檊?�d�$���?       �T�f$@������������������������       �               ��/����?]       ^                    �?      �<       ��#�� @������������������������       �               ��#�� @������������������������       �               z�5��@������������������������       �      ȼ       �cp>@a       f                 �?�r?�L����?       Yk���>)@b       c                  P���?`n����?       � ��w<@������������������������       �               ��#���?d       e                  ���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       /����/#@h       i                  �/�?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ���>��@k       l                     �?`L�Е��?       zVd�t2@������������������������       �               ��/����?m       n                 �Z�?X��qS�?
       �X���0@������������������������       �               0#0#�?������������������������       �      �<	       �P^Cy/@������������������������       �      �       �cp>@q       v                �Y�k�?�w͘�?	       �I����*@r       s                    �?�3`���?       .�r��@������������������������       �               ��#���?t       u                 ����?���`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               �k(��"@x       �                 ?~�?x+2LK�?       ��Z:@@y       �                 ��nZ?z�2|���?       �n�df_7@z       �                 ����?�T�^e��?       =^��:T5@{       �                 }%R?p�BG_��?	       ���M�U3@|                         �Xs?r-�E�T�?       ��<)@}       ~                 p���?h�4���?       �tCP��@������������������������       �               0#0# @������������������������       �               �cp>@�       �                 p�
�?xLU���?       i�ҹ^�@������������������������       �               0����/@�       �                  ���?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?������������������������       �               ���-��@�       �                 p���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                  h��?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?�       �                 p,8�?�����?       ��ȋ_)"@������������������������       �               ��#�� @�       �                 ��B�?X�ih�<�?       ��
@������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?�       �                  ��?�+�bƲ?       =�7*9@�       �                  z��?v=���?       � ��R(@������������������������       �               #0#0&@������������������������       �      ȼ       ��/����?������������������������       �      ��
       ��8��8*@�       �                  �E�?
�f]B�?B       j�Q�>iY@�       �                     �?{|�9�#�?/       zmeGcbQ@�       �                 �8˥?)L垽?       |��[0@������������������������       �        	       ���-��*@�       �                 ��}�?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?�       �                 �Rˡ?ﮃ��y�?$       3�}�J@�       �                 PeT�?!�V���?       <�ٷ0	1@�       �                    �?�֪u�_�?       ��?�8@������������������������       �               0����/@������������������������       �               0#0#�?�       �                 ����?g�wy��?       �f0�v&@������������������������       �               z�5��@�       �                    �?=�N9���?       ��{j�@�       �                 �+tw?      �<       H�4H�4@������������������������       �               0#0#�?������������������������       �               0#0# @�       �                 �C8�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 pt��?vX���<�?       ܐ�VB@�       �                 ����?Jz��܍�?       ۜ�58@�       �                 �S��?xLU���?       ��],7@�       �                 PP��?0�8�4�?       ׁ��t0@�       �                 ���?xLU���?       g�ҹ^�.@�       �                 ͏�?��,���?
       "C�s��,@������������������������       �               /����/#@�       �                 ��U�?���mf�?       寠�?b@�       �                 賆�?v�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �               0#0#�?������������������������       �               ���-��@������������������������       �      �<       ��#���?�       �                   ��?ۼ��?	       �	U�'@�       �                 ���?��n��?       �-H�\@�       �                 �2�o?�֪u�_�?       ��?�8@������������������������       �      ��       0����/@������������������������       �               0#0#�?������������������������       �               ��#���?�       �                 �ߒ�?     ��?       "F�b@������������������������       �               ��#�� @������������������������       �               H�4H�4@�       �                 �=�?���M��?       �Oؽ�@@�       �                 `|W�?���ܤ��?       H4��D6@�       �                  ���?�.�KQu�?       �K̎@������������������������       �               0#0#@������������������������       �               z�5��@������������������������       �        	       �A�A.@�       �                    �?z�G���?       �֔�Э#@�       �                   p��?��[����?       Hl�_A@�       �                 `�k�?�֪u�_�?       ��?�8@�       �                @�~b�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��/���@������������������������       �               0#0#�?������������������������       �               H�4H�4@�       �                 �;�?�I��ҳ�?=       ��s�Y@�       �                 �/��?(d���&�?'       Y%�%�O@�       �                 0��?�Z&s:�?       ~'qγJ@�       �                 ��?jt\���?       �j�O�H@������������������������       �               ��/����?�       �                 �D���|��h�?       �)��%H@�       �                 �~��?�K��t�?       L����"@�       �                 ���?�o���?       o�9�F@������������������������       �               ��#���?������������������������       �               0#0#@�       �                    �?���/��?       V��7�@�       �                  P�"�?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      �<       ��/����?�       �                 `���?��pUз?       ~�w�C@������������������������       �      ȼ       H�4H�48@�       �                 �$/�?��E�B��?	       dߞKC.@������������������������       �               �C=�C=@�       �                 � �?����|e�?       �z �B�@������������������������       �               ��/����?�       �                 0���?X�ih�<�?       ��
@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �      �       �cp>@�       �                ��B�~?%�!�GU�?       m�����%@������������������������       �               ��#�� @�       �                 0ֺ�?�`���6�?       /u��֝!@�       �                 ����?�@G���?       hu��@�       �                    �?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               0����/@������������������������       �               ��#���?�       �                 `G�?      �<       ��+��+D@������������������������       �               H�4H�4@������������������������       �               �z��z�B@�t�b��#     h�hhK ��h��R�(KK�KK��h �B(  �k(��b@��-��bd@�6k�6�c@������a@�+Q��b@�i��R@���b:`@5�@S�X@������C@���b:`@x%jW�vX@�A�A.@��Gp_R@����z�A@        k1��tVQ@�cp>7@        �,����7@��|��,@        ��#�� @���-��@        ��#���?�cp>@        ��#���?                        �cp>@                ��/����?                0����/@        ��#���?��/����?                ��/����?        ��#���?                �k(���5@��/���@        ;��,��@���-��@        ;��,��@��/���@        ��#��@��/����?                ��/����?        ��#��@                ��#���?��/����?                ��/����?        ��#���?                        �cp>@        ��#��0@��/����?                ��/����?        ��#��0@                ^Lg1��F@D�JԮD!@        �#���9@��/����?        ;��,��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        z�5��@                <��,��4@                ���>��,@                z�5��@                ������3@��/���@        ;��,��@��/���@        ��#���?���-��@        ��#���?�cp>@                �cp>@        ��#���?                        ��/���@        ��#��@��/����?        ��#��@                ��#�� @                ��#�� @                        ��/����?        ���>��,@                ��b:��*@                ��#���?                ��#��@��On�(@        ��#���?鰑%@        ��#���?��/����?                ��/����?        ��#���?                        E�JԮD!@        z�5��@��/����?        ��#�� @                ��#���?��/����?        ��#���?                        ��/����?        �>��nK@0����-O@�A�A.@�}�\I@h
��F@��+��+@��k(/D@��]�ڕE@H�4H�4@z�5��@�cp>7@0#0# @z�5��@�cp>7@0#0# @��#�� @/����/3@        ��#���?0����/3@                �cp>'@        ��#���?��/���@        ��#���?                        ��/���@        ��#���?                ��#���?��/���@0#0# @��#���?                        ��/���@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @        �cp>@        z�5��@                Fy�5A@%jW�v%4@0#0#�?Fy�5A@E�JԮD1@0#0#�?�k(��2@��/���.@        <��,��$@��/���.@        ��#�� @0����/@        ��#�� @��/����?                ��/����?        ��#�� @                ��#�� @                z�5��@                        �cp>@        ��#�� @鰑%@        ��#�� @��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                        /����/#@        ��#�� @                ��#���?                ���>��@                �P^Cy/@��/����?0#0#�?        ��/����?        �P^Cy/@        0#0#�?                0#0#�?�P^Cy/@                        �cp>@        ;��,��$@��/����?0#0# @��#���?��/����?0#0# @��#���?                        ��/����?0#0# @        ��/����?                        0#0# @�k(��"@                ��#��@:l��F:2@��+��+$@��#�� @E�JԮD1@0#0#@��#���?E�JԮD1@H�4H�4@        On��O0@H�4H�4@        0����/#@H�4H�4@        �cp>@0#0# @                0#0# @        �cp>@                ���-��@0#0#�?        0����/@                ��/����?0#0#�?        ��/����?                        0#0#�?        ���-��@        ��#���?��/����?                ��/����?        ��#���?                ��#���?        0#0#�?                0#0#�?��#���?                ��#�� @��/����?H�4H�4@��#�� @                        ��/����?H�4H�4@                H�4H�4@        ��/����?                ��/����?H�4H�48@        ��/����?#0#0&@                #0#0&@        ��/����?                        ��8��8*@���>��,@p��F:lI@vb'vb'B@[Lg1��&@
�cp>G@H�4H�4(@        ��/���.@0#0#�?        ���-��*@                ��/����?0#0#�?        ��/����?                        0#0#�?[Lg1��&@��/���>@#0#0&@���>��@�cp>@0#0#@        0����/@0#0#�?        0����/@                        0#0#�?���>��@��/����?H�4H�4@z�5��@                ��#���?��/����?H�4H�4@                H�4H�4@                0#0#�?                0#0# @��#���?��/����?                ��/����?        ��#���?                ��#��@��On�8@�C=�C=@��#���?%jW�v%4@H�4H�4@        %jW�v%4@H�4H�4@        ���-��*@H�4H�4@        ���-��*@0#0# @        ���-��*@0#0#�?        /����/#@                ��/���@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@                        0#0#�?                0#0#�?        ���-��@        ��#���?                z�5��@0����/@0#0#@��#���?0����/@0#0#�?        0����/@0#0#�?        0����/@                        0#0#�?��#���?                ��#�� @        H�4H�4@��#�� @                                H�4H�4@z�5��@0����/@H�4H�48@z�5��@        ��)��)3@z�5��@        0#0#@                0#0#@z�5��@                                �A�A.@        0����/@��+��+@        0����/@0#0# @        0����/@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/���@                        0#0#�?                H�4H�4@z�5��@���-��*@�fm�f�T@z�5��@���-��*@�
��
�E@z�5��@��/���@�ڬ�ڬD@z�5��@0����/@�ڬ�ڬD@        ��/����?        z�5��@��/���@�ڬ�ڬD@z�5��@��/����?0#0#@��#���?        0#0#@��#���?                                0#0#@��#�� @��/����?        ��#�� @��/����?        ��#�� @                        ��/����?                ��/����?                ��/����?�z��z�B@                H�4H�48@        ��/����?��8��8*@                �C=�C=@        ��/����?H�4H�4@        ��/����?                ��/����?H�4H�4@        ��/����?                        H�4H�4@        �cp>@        z�5��@�cp>@0#0# @��#�� @                ��#���?�cp>@0#0# @        �cp>@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @        0����/@        ��#���?                                ��+��+D@                H�4H�4@                �z��z�B@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ� �thFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK߅�h��B�0         T                 �j"�?J��r�D�?)      c?���m}@       E                 p��?�R�d�?l       # mnf@       B                  �h?�� Բ�?X       �c��Na@       ?                 `ٯ�?>��5s��?S       ��(-`@       $                  �g<�?�M�����?O       	i!o^@       !                 ���G?�օ����?'       8��%ǦM@                        ���s?���/��?       �JX���F@                        ��IL?��f�n�?       5(q�GA@	       
                  `���?�_�A�?       肵�e`@������������������������       �               ��/����?������������������������       �               ;��,��@                        0a?��|��?       ���ĺw;@������������������������       �               ��/���@                        �*%?l%@�"�?       ��[�7@                        �1?,��c`�?       &��t5)@������������������������       �               鰑%@                        �!"?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?                        ���u?4k�"O��?       �?<��*&@������������������������       �               z�5��@                        �[�Z?, k�Lj�?       �q��l}@������������������������       �               �cp>@                        �p�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?                            �?����X��?	       &��֞&@                         `�J�?~d�$���?       �T�f@                        �؉�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       z�5��@������������������������       �               z�5��@"       #                    �?      �<       ���-��*@������������������������       �               ��On�(@������������������������       �               ��/����?%       (                 @I��>�FL�?�?(       OO�{7O@&       '                 �#�>jQ��?       �s�=�!@������������������������       �               ��#�� @������������������������       �               ���-��@)       4                    �?4D@�%�?!       2Wd��J@*       +                  �~��?� ��i�?       �u�:hA@������������������������       �               ��/����?,       -                 �:W>?L�7Ke��?       �B�n�@@������������������������       �      ��       
�#���9@.       3                 ���?���/��?       U��7�@/       2                 ؽkz?�d�$���?       �T�f@0       1                 �
<P?      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@������������������������       �      ȼ       ��/����?������������������������       �               �cp>@5       <                 �/?�KĈ�?       y�Zc�2@6       7                 �?�)z� ��?	       ��\�,@������������������������       �               z�5��@8       ;                 'uk?Δfm���?       ��Z�N@9       :                 Ш��?�`@s'��?       Ei_y,*@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               ��#���?=       >                  ��?      �<       0����/@������������������������       �               ��/����?������������������������       �               ��/���@@       A                    �?      �<       ��/���@������������������������       �               �cp>@������������������������       �               0����/@C       D                  �.�?�*�'=P�?        �2"@������������������������       �               0#0# @������������������������       �      ȼ       ��/����?F       M                 ���x?
��ɝO�?       p�� ��D@G       L                 0A��?��2eK�?	       <=h��.@H       I                 远�?p��H��?       v�I�@������������������������       �               �cp>@J       K                 �2OF?����?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?������������������������       �               0#0# @N       S                 �-��?���~�Q�?       A���6 :@O       R                   E(�? LD1�ӳ?
       ����8@P       Q                 �ا�?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �               鰑5@������������������������       �               0#0#�?U       �                 �LW�?�Qr����?�       ^/)?O6r@V                         `���?�a�&���?B       �#�[@W       `                  �mS?��o��C�?,       T��^HVR@X       Y                  ;��?���+���?       ��=��'@������������������������       �               z�5��@Z       _                 ТO?P�H�q�?       ��	0�!@[       \                 h꟫?��n��?       �-H�\@������������������������       �               0����/@]       ^                 ����?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               0#0# @a       |                  �?�hd��z�?&       �~�U�N@b       c                 0=T�?�W�w��?#       y;���K@������������������������       �               0#0#�?d       e                 �vs?�����?"       a���"K@������������������������       �        	       �P^Cy/@f       w                 p)�w?�~"�4�?       ��⃃_C@g       t                 �#��?���'>y�?       Y0ӝ�*4@h       k                 �Z�?xR�wrA�?       w���&J1@i       j                 ��v�?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?l       m                  p���?�b���:�?
       �
#���,@������������������������       �               ��/����?n       s                 hU�<?*PThD]�?	       �p�]�*@o       p                 @�A�?�f@���?       hy���"@������������������������       �      ȼ       z�5��@q       r                ����?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               ��#��@u       v                 �vQ?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?x       {                 �g\�?�wV����?       Bi�i�2@y       z                 �t�?�f@���?       hy���"@������������������������       �      ��       ���>��@������������������������       �               0#0# @������������������������       �               �k(��"@}       ~                 P�`�?�D#���?       �B�j@������������������������       �               0#0#@������������������������       �               ��#�� @�       �                    �?0�a(I��?       T�>��wB@�       �                  ��a?DUK&�?       $I/���<@�       �                 ���?����?       �g=�2@�       �                 �Z�?�yoJ	�?       ���8
�0@�       �                   Y��?�)��R=�?       �
3�e1)@�       �                  �0��?��n��?       �-H�\@�       �                ��?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �               0����/@������������������������       �               ��#���?�       �                 pG˘?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/���@�       �                 �;��?�J���?       ��*]Y@������������������������       �               ��#�� @������������������������       �               0#0# @������������������������       �      �<       ��#�� @������������������������       �               ��+��+$@�       �                 ����?a�ox��?       
c��0 @������������������������       �               ��#���?�       �                 X��?      �<       �C=�C=@������������������������       �               0#0# @������������������������       �               ��+��+@�       �                 �%r�?���JeF�?{       9ϊl��f@�       �                 P�ʏ?N�o$���?\       ����\a@�       �                 ��{�?�v����?%       �H<OB�I@������������������������       �               ��+��+@�       �                 `���?�,����?!       �ж��rG@�       �                 ���? ��k~�?       X�3Á�E@�       �                 ����?������?       ǈ��&mB@�       �                  �@�?��7^�6�?       �IU��=@������������������������       �               ��#���?�       �                 �5�z?��, �#�?       ��
���<@������������������������       �               ��#���?�       �                  -��?�R�Gz۱?       ��P��;@������������������������       �               ���-��:@������������������������       �               0#0#�?�       �                  �JV�?�Qk��?       ��Th!�@������������������������       �               ��/����?�       �                 ��λ?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?�       �                ����}?�)z� ��?       �\�@�       �                    �?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �      м       ��/����?�       �                 ����?      �<       H�4H�4@������������������������       �               0#0#�?������������������������       �               0#0# @�       �                 �6SZ?l�}����?7       ��h��U@�       �                  ���?�H�F��?       J2�$��D@�       �                 `;ĝ?v�GZ��?       N+A2?@������������������������       �               ��/���@�       �                 px��?H��aB��?       y/�t�/;@�       �                 `�v�?���zc�?       1��.D+9@�       �                 0"��?W�|!��?       \�pq�T5@�       �                  ��?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@�       �                 `(¢?�x�<�?	       X&b��q1@������������������������       �               ZLg1��&@�       �                 $��?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#��@�       �                 h�I�?      �<       ��/���@������������������������       �               ��/����?������������������������       �               �cp>@������������������������       �               0#0# @�       �                 �`��?�}/W�?       �r�.�%@�       �                 PeT�?��^���?       ���w!@������������������������       �               0#0# @������������������������       �      ��       ���-��@������������������������       �               0#0# @�       �                 p�:�?_����?       ��_�
�F@�       �                 ��?|��`p��?	       �����'@�       �                  ��?l*�'=P�?        �2"@������������������������       �               �C=�C=@�       �                    �?x�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �      ȼ       �cp>@������������������������       �      ��       B�A�@@�       �                   �0�? ��ճC�?       鰑E@�       �                 @�%�?���};��?	       ��;̑�%@������������������������       �               ��/����?�       �                 ��?d*�'=P�?        �2"@������������������������       �               H�4H�4@�       �                8�fG�?z��`p��?       �����@������������������������       �               0#0#�?�       �                 @8��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 �&��?      �<       =�C=�C?@������������������������       �               0#0# @������������������������       �               �s?�s?=@�t�bh�hhK ��h��R�(KK�KK��h �B�  �YLg1b@t�H���e@�LɔL	c@"�}��P@�h
�W@vb'vb'2@���b:P@���|�P@0#0# @���b:P@Pn��OP@        ���b:P@��|��L@        �,����7@����z�A@        �,����7@h
��6@        ��b:��*@鰑5@        ;��,��@��/����?                ��/����?        ;��,��@                ��#�� @/����/3@                ��/���@        ��#�� @��/���.@        ��#���?�cp>'@                鰑%@        ��#���?��/����?        ��#���?                        ��/����?        ���>��@��/���@        z�5��@                ��#���?��/���@                �cp>@        ��#���?��/����?                ��/����?        ��#���?                <��,��$@��/����?        ��#��@��/����?        ��#���?��/����?                ��/����?        ��#���?                z�5��@                z�5��@                        ���-��*@                ��On�(@                ��/����?        ��k(/D@h
��6@        ��#�� @���-��@        ��#�� @                        ���-��@        d:��,&C@��/���.@        Jp�}>@0����/@                ��/����?        Kp�}>@��/���@        
�#���9@                ��#��@��/���@        ��#��@��/����?        ��#��@                ��#���?                z�5��@                        ��/����?                �cp>@        ��#�� @鰑%@        ��#�� @�cp>@        z�5��@                ��#�� @�cp>@        ��#���?�cp>@                �cp>@        ��#���?                ��#���?                        0����/@                ��/����?                ��/���@                ��/���@                �cp>@                0����/@                ��/����?0#0# @                0#0# @        ��/����?        z�5��@�a#6�;@��+��+$@z�5��@��/���@0#0# @z�5��@��/���@                �cp>@        z�5��@��/����?        z�5��@                        ��/����?                        0#0# @        �e�_��7@0#0# @        �e�_��7@0#0#�?        �cp>@0#0#�?        �cp>@                        0#0#�?        鰑5@                        0#0#�?���khS@h
���S@K`F`�`@.�����K@鰑5@B�A�@@|�5��H@鰑%@��8��8*@��#��@0����/@H�4H�4@z�5��@                ��#���?0����/@H�4H�4@��#���?0����/@0#0#�?        0����/@        ��#���?        0#0#�?��#���?                                0#0#�?                0#0# @]Lg1��F@�cp>@��+��+$@�k(���E@�cp>@H�4H�4@                0#0#�?�k(���E@�cp>@��+��+@�P^Cy/@                *�����;@�cp>@��+��+@ZLg1��&@�cp>@H�4H�4@[Lg1��&@�cp>@H�4H�4@        ��/����?0#0#�?        ��/����?                        0#0#�?ZLg1��&@��/����?0#0# @        ��/����?        [Lg1��&@        0#0# @���>��@        0#0# @z�5��@                ��#���?        0#0# @��#���?                                0#0# @��#��@                        �cp>@                ��/����?                ��/����?        ��#��0@        0#0# @���>��@        0#0# @���>��@                                0#0# @�k(��"@                ��#�� @        0#0#@                0#0#@��#�� @                z�5��@鰑%@��+��+4@;��,��@鰑%@��8��8*@;��,��@鰑%@H�4H�4@z�5��@鰑%@H�4H�4@��#���?鰑%@0#0#�?��#���?0����/@0#0#�?        0����/@0#0#�?                0#0#�?        0����/@        ��#���?                        �cp>@                ��/����?                ��/���@        ��#�� @        0#0# @��#�� @                                0#0# @��#�� @                                ��+��+$@��#���?        �C=�C=@��#���?                                �C=�C=@                0#0# @                ��+��+@�k(���5@H�)�BM@p�6k�6Y@�k(���5@�a#6�K@.��+��N@z�5��@On��O@@��8��8*@                ��+��+@z�5��@Pn��O@@0#0# @z�5��@On��O@@��+��+@��#�� @�_��e�=@��+��+@��#�� @���-��:@0#0#�?��#���?                ��#���?���-��:@0#0#�?��#���?                        ���-��:@0#0#�?        ���-��:@                        0#0#�?        �cp>@0#0#@        ��/����?                ��/����?0#0#@                0#0#@        ��/����?        ��#��@�cp>@        ��#��@��/����?        ��#��@                        ��/����?                ��/����?                        H�4H�4@                0#0#�?                0#0# @�P^Cy/@�cp>7@J�4H�4H@�P^Cy/@/����/3@�C=�C=@�P^Cy/@��On�(@H�4H�4@        ��/���@        �P^Cy/@E�JԮD!@H�4H�4@�P^Cy/@D�JԮD!@0#0#�?�P^Cy/@0����/@0#0#�?        �cp>@0#0#�?                0#0#�?        �cp>@        �P^Cy/@��/����?        ZLg1��&@                ��#��@��/����?                ��/����?        ��#��@                        ��/���@                ��/����?                �cp>@                        0#0# @        ���-��@0#0#@        ���-��@0#0# @                0#0# @        ���-��@                        0#0# @        ��/���@�ڬ�ڬD@        ��/���@0#0# @        ��/����?0#0# @                �C=�C=@        ��/����?0#0#�?                0#0#�?        ��/����?                �cp>@                        B�A�@@        �cp>@������C@        �cp>@0#0# @        ��/����?                ��/����?0#0# @                H�4H�4@        ��/����?0#0# @                0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?                =�C=�C?@                0#0# @                �s?�s?=@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��1hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKم�h��Bx/         |                  ��d�?#�q�>�?%      X�y�l}@       _                 �4�?vP�հ��?�       p����8k@       F                 ��U�?��ױ��?u       M�eZf@                        `�]?�H����?[       6��[�a@                        ��?#����?       v�߄�3@                        ��x?��t� �?       ����x&@                         �P��?�FO���?       �ߌ$@������������������������       �               ;��,��@	       
                  �g<�?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �               ��#�� @       E                 @�˒?��& ��?P       ���n��^@                        �$I�?#�@���?I       ���˴[@������������������������       �               ���>��@       :                 ��r?��q�C�?F       ����Y@       9                 p���?���/x��?9       ���l��T@       $                 ����?P�w3���?6       �N
��S@       #                 ��$�?�H�����?       K��XE@                        @F��~q����?       �w��D@                        ��j?P���i�?       �#���=@                           �?�`���6�?       .u��֝!@                       @� 4$?�`@s'��?       Ei_y,*@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               0#0# @                         �A?      �<       鰑5@������������������������       �               ��/���@������������������������       �               D�JԮD1@                         ���T?Ԕfm���?       �0��z'@������������������������       �               z�5��@!       "                 Pkf?      �<       D�JԮD!@������������������������       �               ��/���@������������������������       �               0����/@������������������������       �      �<       ��#���?%       6                   �P�?J��`�?       z�_P�A@&       3                 �q�3?8>Í�`�?       &��3�Q>@'       (                 ���x?b�N�?       �Ȓ���2@������������������������       �               ;��,��@)       0                 ��Yk?����p��?
       �˰�\C+@*       -                 h�ف?�n�l���?       ���5F'@+       ,                 �e?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?.       /                  ��?x5JH���?       �MOI#@������������������������       �               E�JԮD!@������������������������       �               0#0#�?1       2                 ��-�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?4       5                 p�37?      �<	       �cp>'@������������������������       �               ��/����?������������������������       �               鰑%@7       8                 \F�M?      �<       ;��,��@������������������������       �               z�5��@������������������������       �               ��#�� @������������������������       �               ;��,��@;       B                 �p�U?�>Kn$P�?       1�L\�84@<       ?                 PFsf?��{@��?       ��I�@2@=       >                 ��\�?$ k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?@       A                 �4C�?h�s�	�?       f���*@������������������������       �      �<       z�5��(@������������������������       �      ȼ       ��/����?C       D                 v� �?��G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               {�5��(@G       \                 0�ݮ?N0��S�?       qӵ�%B@H       K                  �9��?i�z��P�?       ?0F��m;@I       J                 ���?�}	;	�?       uK�>4%@������������������������       �      ��       0����/#@������������������������       �               0#0#�?L       W                 ��U�?��ҭ�x�?       �
�H��0@M       T                 p��?�]
���?	       ��Ј�'@N       O                 �CǨ?~�G���?       '5L�`�@������������������������       �               0#0# @P       Q                 py��?�@G���?       hu��@������������������������       �               ��/����?R       S                 n�h?z�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?U       V                 ��?�D�-,�?       �D'ŰO@������������������������       �               ��#���?������������������������       �               ��+��+@X       [                 @?���mf�?       毠�?b@Y       Z                 n(�?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �               ��/����?]       ^                 �j��?      �<       D�JԮD!@������������������������       �               ��/����?������������������������       �               ���-��@`       e                   ���?��7�Jt�?       x�@��yC@a       d                 @��?��^���?       ���w!@b       c                 x�P�?      �<       ���-��@������������������������       �               ��/����?������������������������       �               �cp>@������������������������       �               0#0# @f       {                 @���?$ȇ��?       ��8>@g       n                 (D�?���v� �?       p���3@h       i                    �?&�b���?       �GXvƒ@������������������������       �               ��/����?j       m                 ��x�?��ڰ�x�?       �K�f�@k       l                 `'v�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               ��#��@o       z                  ����?�]
���?
       ��Ј�'@p       q                 �@�?���3�?	       &��X&@������������������������       �               ��/����?r       y                 �V"P?޾�R���?       :�S) $@s       t                 0V�?:�N9���?       ��{j�@������������������������       �               ��/����?u       x                  ���?b,���O�?       ���/>@v       w                      �J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               0#0# @������������������������       �               ��+��+@������������������������       �      м       ��/����?������������������������       �               #0#0&@}       �                 ���?�\��
�?�       R�h�o@~       �                 �y���#��e��?)       �� �~Q@       �                 8r�t?|+�r7��?       ؖ��<5@@�       �                  L��?��$�<�?       P���4:@�       �                 �+>\?l��H��?       v�I�@������������������������       �               ��/���@������������������������       �      �<       z�5��@�       �                   ��?�� N��?	       �L�EBC3@������������������������       �               ��/���.@�       �                 �<�l?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@�       �                 ��=�?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ;��,��@�       �                 �f�V?v�xrI��?       �RFu!�B@�       �                ���?�N,u��?       ��u�=@�       �                  2��?DBms�?       ��֖��;@�       �                 p|�}?�q�Ptܳ?       Q�� 5�7@������������������������       �               ��b:��*@�       �                 ��q�?�FO���?       �ߌ$@������������������������       �               �k(��"@������������������������       �      ȼ       ��/����?�       �                 � ��?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@������������������������       �      ȼ       ��/����?�       �                 pU�\?���`�?       ��
�Me@������������������������       �               0����/@�       �                 ��Y�?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?�       �                   �0�?��5\�9�?l       ���f@�       �                 �T�Z?z���6�?       Q��a�DH@�       �                 @�=�?H���@�?       �CA�9[;@�       �                 �D��?�zœ���?       HG���t0@������������������������       �               0#0#@������������������������       �      м       z�5��(@�       �                 CJ�?f�/W�D�?       ���z^�%@������������������������       �               0#0#@�       �                 ����?��|��?       ���ĺw@������������������������       �               ��#���?�       �                 @�ſ?l@ȱ��?       om���S@������������������������       �               0����/@������������������������       �               ��#���?������������������������       �      Լ       ��-��-5@�       �                 ���?���7RN�?S       $�^{��`@�       �                   Y��?ܙ�X�t�?%       �#�O@�       �                 @Ws�?������?       2�<��@@�       �                 `bp�?d����?       �����!@������������������������       �               ��/����?������������������������       �      ��       �C=�C=@�       �                 ��?�^����?       �y���!8@�       �                 R{�?����*�?
       �	�c/(+@�       �                ���?�}	;	�?       uK�>4%@������������������������       �               /����/#@������������������������       �               0#0#�?�       �                 p�
�?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               鰑%@�       �                 pyXE?�3"�b��?       ���w�<@�       �                  @�a�?\������?       ��Iē'@�       �                ���u?`%��̫�?       �@�o#@�       �                 �+.�?�;[��G�?       �O�;�]!@������������������������       �      ��       ���-��@�       �                  0p��?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ܼ       ��#���?������������������������       �               ��#�� @������������������������       �      ��       S2%S2%1@�       �                 @� ?�aM��t�?.       5�2�	R@�       �                 ȯ�?��jN�?       >@
�>@������������������������       �               ��/����?�       �                ����?�nl4�/�?       SBe+�1<@�       �                 �"�?�s�R�͵?       �o�97@�       �                 ����?�o���?       o�9�F@������������������������       �               0#0#@������������������������       �               ��#���?������������������������       �               vb'vb'2@�       �                  L��?��`i��?       �؛.�@�       �                 �ec�?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               0#0# @�       �                 �^��?Pp	�/��?       J�YŦ'E@�       �                    �?      �<       =�C=�C?@������������������������       �        	       �A�A.@������������������������       �        
       0#0#0@�       �                 ����?�^�F�M�?       ��ޚ�&@������������������������       �               ��/����?������������������������       �               ��+��+$@�t�bh�hhK ��h��R�(KK�KK��h �BX  YUUUU5a@�xr�'we@��+��+d@��k(/T@�D�J�.Y@xb'vb'B@�k(��R@�'�xr�V@�C=�C=,@��Gp_R@Qn��OP@0#0#@��,���1@��/����?        �k(��"@��/����?        �k(��"@��/����?        ;��,��@                ��#��@��/����?                ��/����?        ��#��@                        ��/����?        ��#�� @                -�����K@�]�ڕ�O@0#0#@�k(���E@�]�ڕ�O@0#0#@���>��@                �YLg1B@�]�ڕ�O@0#0#@\Lg1��6@��|��L@H�4H�4@��,���1@��|��L@H�4H�4@;��,��@����z�A@0#0# @��#��@����z�A@0#0# @��#���?���-��:@0#0# @��#���?�cp>@0#0# @��#���?�cp>@        ��#���?                        �cp>@                        0#0# @        鰑5@                ��/���@                D�JԮD1@        z�5��@D�JԮD!@        z�5��@                        D�JԮD!@                ��/���@                0����/@        ��#���?                |�5��(@h
��6@0#0#�?���>��@h
��6@0#0#�?���>��@鰑%@0#0#�?;��,��@                ��#�� @鰑%@0#0#�?��#���?0����/#@0#0#�?��#���?��/����?        ��#���?                        ��/����?                D�JԮD!@0#0#�?        E�JԮD!@                        0#0#�?��#���?��/����?                ��/����?        ��#���?                        �cp>'@                ��/����?                鰑%@        ;��,��@                z�5��@                ��#�� @                ;��,��@                ��b:��*@�cp>@0#0#�?��b:��*@0����/@        ��#���?��/���@                ��/���@        ��#���?                z�5��(@��/����?        z�5��(@                        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?{�5��(@                ��#���?��On�8@��+��+$@��#���?On��O0@��+��+$@        0����/#@0#0#�?        0����/#@                        0#0#�?��#���?���-��@vb'vb'"@��#���?�cp>@0#0# @        �cp>@H�4H�4@                0#0# @        �cp>@0#0#�?        ��/����?                ��/����?0#0#�?                0#0#�?        ��/����?        ��#���?        ��+��+@��#���?                                ��+��+@        ��/���@0#0#�?        �cp>@0#0#�?                0#0#�?        �cp>@                ��/����?                D�JԮD!@                ��/����?                ���-��@        z�5��@鰑%@#0#06@        ���-��@0#0# @        ���-��@                ��/����?                �cp>@                        0#0# @z�5��@��/���@��+��+4@z�5��@��/���@vb'vb'"@;��,��@��/����?0#0#�?        ��/����?        ;��,��@        0#0#�?��#���?        0#0#�?��#���?                                0#0#�?��#��@                ��#���?�cp>@0#0# @��#���?��/����?0#0# @        ��/����?        ��#���?��/����?0#0# @��#���?��/����?H�4H�4@        ��/����?        ��#���?        H�4H�4@��#���?        0#0#�?��#���?                                0#0#�?                0#0# @                ��+��+@        ��/����?                        #0#0&@v�}wL@¬��z�Q@C�C=�C_@�k(��B@��/���>@0#0# @<��,��$@h
��6@        ��#��@h
��6@        z�5��@��/���@                ��/���@        z�5��@                ��#���?:l��F:2@                ��/���.@        ��#���?�cp>@        ��#���?                        �cp>@        z�5��@                ��#���?                ;��,��@                ��b:��:@E�JԮD!@0#0# @�#���9@��/���@        �#���9@��/����?        [Lg1��6@��/����?        ��b:��*@                �k(��"@��/����?        �k(��"@                        ��/����?        z�5��@��/����?                ��/����?        z�5��@                        ��/����?        ��#���?0����/@0#0# @        0����/@        ��#���?        0#0# @                0#0# @��#���?                ������3@'jW�v%D@2��+��^@���>��,@0����/@�s?�s?=@���>��,@0����/@0#0# @{�5��(@        0#0#@                0#0#@z�5��(@                ��#�� @0����/@0#0#@                0#0#@��#�� @0����/@        ��#���?                ��#���?0����/@                0����/@        ��#���?                                ��-��-5@;��,��@����z�A@2��-�rW@z�5��@��/���>@�C=�C=<@        �cp>7@��+��+$@        ��/����?�C=�C=@        ��/����?                        �C=�C=@        鰑5@H�4H�4@        鰑%@H�4H�4@        /����/#@0#0#�?        /����/#@                        0#0#�?        ��/����?0#0# @        ��/����?                        0#0# @        鰑%@        z�5��@��/���@vb'vb'2@z�5��@��/���@0#0#�?��#���?��/���@0#0#�?        ��/���@0#0#�?        ���-��@                ��/����?0#0#�?        ��/����?                        0#0#�?��#���?                ��#�� @                                S2%S2%1@��#�� @0����/@9��8�cP@��#�� @��/���@H�4H�48@        ��/����?        ��#�� @��/����?H�4H�48@��#���?        #0#06@��#���?        0#0#@                0#0#@��#���?                                vb'vb'2@��#���?��/����?0#0# @��#���?��/����?        ��#���?                        ��/����?                        0#0# @        ��/����?�ڬ�ڬD@                =�C=�C?@                �A�A.@                0#0#0@        ��/����?��+��+$@        ��/����?                        ��+��+$@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�JIhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKم�h��Bx/         �                 `r�t?��8�@�?)      ;�ZH��}@       �                 ��C?6�ǥ#p�?�       ��jxhv@       n                   �0�?Rs��w"�?�       ��?�q@       W                  4�?\��k<�?~       �]2l�.h@       B                 @�ő?�i5�gS�?b       �I���c@       9                 0�,7?�e΅��?N       /DP��^@       8                  �_�?�Р�k��?D       ,�Y@       +                 ~`�����1��?;       =�ߋ2V@	                        �$?Z?��g���?$       #C.�yH@
                        0��\?��k*���?       ���b-@                         �.�?���3�?       ���(+�%@                        ���`?r@ȱ��?       om���S@������������������������       �               0����/@������������������������       �               ��#���?                        �N�L?ޗZ�	7�?       j~���@������������������������       �               z�5��@������������������������       �      �<       ��/����?������������������������       �               ��/���@                          �G�?
<4BL��?       �G.�� A@                        ��?l@ȱ��?       nm���S@������������������������       �               ��#���?������������������������       �      ��       0����/@       &                 `�j�?b�6P$g�?       4^��l<@                        �<��>��x_F-�?       x%jW�v8@������������������������       �               ��/����?       %                  ��?XՏ�m|�?       ��h
�7@       "                 �@�?��E�B��?       �'�xr�6@                        ���|?k� ѽ?	       �����.@������������������������       �               <��,��$@                           �?~d�$���?       �T�f@������������������������       �               ��#���?        !                  ���?����?       ��X�)B@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?#       $                 Z��?�_�A�?       肵�e`@������������������������       �               ��/����?������������������������       �               ;��,��@������������������������       �      �<       ��/����?'       (                 p���?J��NV=�?       �t�ܲ@������������������������       �               0#0#�?)       *                �J��?f%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?,       -                 ���	?�s���?       ZE��K�C@������������������������       �               ��b:��*@.       5                 pt$x?^(��I�?       d#6�a:@/       0                 ���X?`����?       �Fx�v�5@������������������������       �               ��/����?1       4                �н��?�FO���?       �ߌ4@2       3                 `Qd�>      �<
       �k(��2@������������������������       �               ��#���?������������������������       �        	       ��,���1@������������������������       �      ȼ       ��/����?6       7                 X���?6 k�Lj�?       �q��l}@������������������������       �      �<       ��/���@������������������������       �               ��#���?������������������������       �        	       ��b:��*@:       A                 p��A?Nͻ�&��?
       |���g�1@;       <                 ���g?tf�T6|�?       x,*��P+@������������������������       �               �cp>@=       @                 @F�8ǵ3���?       �q�ͨ�@>       ?                 q� ?��|��?       ���ĺw@������������������������       �               ��#�� @������������������������       �               0����/@������������������������       �               ��#���?������������������������       �               ��#��@C       D                 @�#�?����lB�?       ,��	�hB@������������������������       �               0#0#@E       V                 `3L�?dv��&�?       �=�Ìd@@F       U                 ���@?�ls���?       ��2�Ax7@G       H                 �A��?^r�.���?       x6.��s5@������������������������       �               ��/����?I       N                 �ѓ?���v���?       ��ԽI~4@J       K                 �U�?�d�$���?       �T�f@������������������������       �               ��#�� @L       M                 `U�?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?O       R                  �P��?X����1�?
       �l����.@P       Q                  p%+�?      �<       �k(��"@������������������������       �               ��#���?������������������������       �               ��#�� @S       T                 ����?�D�-,�?       �D'ŰO@������������������������       �               ��#���?������������������������       �               ��+��+@������������������������       �               0#0# @������������������������       �      ȼ       �k(��"@X       e                 Pz9�?D3�h���?       6QpԂKB@Y       Z                 ����?Ի�$�+�?       v��;k4@������������������������       �               0#0# @[       \                 _%?2N���?       /0۽�f2@������������������������       �      ��
       ���-��*@]       `                 �U�<?��`i��?       �؛.�@^       _                 @��8?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?a       b                    �?�� ��?       rp� k@������������������������       �               ��/����?c       d                 p��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?f       k                 �$|�?H�b̒0�?       ���+0@g       h                  PV��?U
�6���?       Z�4�#R"@������������������������       �               ;��,��@i       j                 ��?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@l       m                 ���?d�ih�<�?       ��
@������������������������       �               ��/����?������������������������       �               H�4H�4@o       �                 S1�?+F���?2       ���%�S@p       �                    �?0ƞ���?$       U^s��I@q       �                 ��h�?�o�·<�?       �&�g?@r       }                 ��N�?�)z� ��?       ��\�<@s       |                 �;̑?�����?       ��/̸I3@t       {                 @?^n����?       Ԁh��K.@u       z                  t�޾�_�A�?       肵�e`,@v       w                 �e�O?���/��?       V��7�@������������������������       �               �cp>@x       y                 �`3x?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �               z�5��@������������������������       �      м       ��/����?������������������������       �               ��#��@~       �                  �`<?vQ��?       �s�=�!@       �                  `<��?h�r{��?       e�6� @�       �                 ��	r?      �<       0����/@������������������������       �               ��/����?������������������������       �               ��/���@�       �                 �M��?b%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �               H�4H�4@�       �                 ����?x�1q�X�?       ���!�4@�       �                 ����?:4|���?       	�T|qt2@�       �                 ���?��I@�?	       �2d�%@�       �                 Yu?�(���?       y��uk!@������������������������       �               ��#���?������������������������       �               ��/���@�       �                 P[��?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?������������������������       �      ��       ��/���@�       �                  �E�?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?�       �                    �?      �<       �;�;;@������������������������       �               H�4H�4(@������������������������       �        	       �A�A.@�       �                  ��?�z�R�?5       =�[�؏U@�       �                  1�?����BW�?,       �]�J�Q@�       �                 ��j�?�G�N�J�?       jX\�=@�       �                 �@�?X�ђ���?       �oFݜh5@������������������������       �               ��/���@�       �                  `��?��|��?       ���ĺw+@������������������������       �               ��#�� @�       �                 @F�p@ȱ��?
       om���S'@�       �                  ���?Δfm���?       ��Z�N@�       �                 �fQ?�`@s'��?       Ei_y,*@������������������������       �               �cp>@�       �                 p'v�?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               ��#���?������������������������       �               ��/���@�       �                 ����?��6L�n�?       �E#��h @�       �                 `�??�d�$���?       �T�f@������������������������       �               ��#�� @�       �                ��+��?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               z�5��@�       �                 0��?�J�>��?       .��
RD@�       �                 p�~t?&�g���?       ��u3@�       �                  ��`?b,���O�?       ���/>@������������������������       �               ��#���?������������������������       �               H�4H�4@�       �                 0�"]?����VV�?	       A�R.�.@������������������������       �      �<       ��|��,@������������������������       �               0#0#�?�       �                 @�Q?�G�,.̷?       �J�$r.5@�       �                 �U*P?)���?       y��uk!@������������������������       �               ��/���@������������������������       �               ��#���?�       �                 �.KR?      �<       ��On�(@������������������������       �               ��/����?������������������������       �               �cp>'@�       �                 ��Z�?X�4X��?	       �<�?p�/@�       �                  y��?�\z����?       ���U��!@�       �                 0�
�?�w��d��?       �0���s@�       �                ���(z?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               �cp>@������������������������       �               ��#�� @������������������������       �               �C=�C=@�       �                 �6Sz?H���h!�?D       �m�u�d\@�       �                   ��?*^�yU�?       ��7�1�#@������������������������       �               ��/����?�       �                  �~��?w�;B��?       ՟���	 @������������������������       �               ��+��+@�       �                  ���?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 p6��?@)�虶?>       z�D��Y@������������������������       �      ȼ%       �C=�C=L@�       �                 �|�?l�Ld�?       F����G@������������������������       �               �cp>@�       �                  ��d�?�~���9�?       �q�Ί#F@�       �                 @��?|��`p��?       �����@�       �                 �1��?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               H�4H�4@������������������������       �      ȼ       ��)��)C@�t�bh�hhK ��h��R�(KK�KK��h �BX  �5��P>b@�+Q��b@�����f@�5��P>b@����z�a@gJ�dJ�Q@�P^CyM`@�H��tXU@�C=�C=L@�>��n[@H�)�BM@k�6k�69@�#���Y@�)�B�D@H�4H�4(@�b:���S@������C@0#0#�?�YLg1R@��|��<@0#0#�?    �M@��|��<@0#0#�?�#���9@h
��6@0#0#�?��#��@鰑%@        ��#��@���-��@        ��#���?0����/@                0����/@        ��#���?                z�5��@��/����?        z�5��@                        ��/����?                ��/���@        �k(���5@�cp>'@0#0#�?��#���?0����/@        ��#���?                        0����/@        <��,��4@���-��@0#0#�?������3@0����/@                ��/����?        ������3@��/���@        ������3@�cp>@        ���>��,@��/����?        <��,��$@                ��#��@��/����?        ��#���?                z�5��@��/����?        z�5��@                        ��/����?        ;��,��@��/����?                ��/����?        ;��,��@                        ��/����?        ��#���?��/����?0#0#�?                0#0#�?��#���?��/����?                ��/����?        ��#���?                ��#��@@���-��@        ��b:��*@                ������3@���-��@        �k(��2@�cp>@                ��/����?        �k(��2@��/����?        �k(��2@                ��#���?                ��,���1@                        ��/����?        ��#���?��/���@                ��/���@        ��#���?                ��b:��*@                ���>��@鰑%@        z�5��@鰑%@                �cp>@        z�5��@0����/@        ��#�� @0����/@        ��#�� @                        0����/@        ��#���?                ��#��@                �,����7@��/����?#0#0&@                0#0#@�,����7@��/����?�C=�C=@���>��,@��/����?�C=�C=@���>��,@��/����?��+��+@        ��/����?        ���>��,@��/����?��+��+@��#��@��/����?        ��#�� @                ��#�� @��/����?        ��#�� @                        ��/����?        ;��,��$@        ��+��+@�k(��"@                ��#���?                ��#�� @                ��#���?        ��+��+@��#���?                                ��+��+@                0#0# @�k(��"@                z�5��@E�JԮD1@��8��8*@��#���?��/���.@0#0#@                0#0# @��#���?��/���.@0#0# @        ���-��*@        ��#���?��/����?0#0# @��#���?        0#0#�?                0#0#�?��#���?                        ��/����?0#0#�?        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?;��,��@��/����?vb'vb'"@;��,��@��/����?H�4H�4@;��,��@                        ��/����?H�4H�4@        ��/����?                        H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@<��,��4@���-��:@=�C=�C?@=��,��4@���-��:@0#0#@��#��0@�cp>'@H�4H�4@��#��0@�cp>'@        ���>��,@0����/@        <��,��$@0����/@        <��,��$@��/���@        ��#��@��/���@                �cp>@        ��#��@��/����?        ��#��@                        ��/����?        z�5��@                        ��/����?        ��#��@                ��#�� @���-��@        ��#���?���-��@                0����/@                ��/����?                ��/���@        ��#���?��/����?        ��#���?                        ��/����?        ��#���?                                H�4H�4@��#��@��/���.@0#0#�?z�5��@��/���.@        z�5��@��/���@        ��#���?��/���@        ��#���?                        ��/���@        ��#�� @                ��#���?                ��#���?                        ��/���@        ��#���?        0#0#�?                0#0#�?��#���?                                �;�;;@                H�4H�4(@                �A�A.@�P^Cy/@M!�ML@�C=�C=,@��b:��*@c#6�aJ@0#0#@ZLg1��&@:l��F:2@        ��#��@E�JԮD1@                ��/���@        ��#��@/����/#@        ��#�� @                ��#�� @/����/#@        ��#�� @�cp>@        ��#���?�cp>@                �cp>@        ��#���?�cp>@                �cp>@        ��#���?                ��#���?                        ��/���@        ���>��@��/����?        ��#��@��/����?        ��#�� @                ��#�� @��/����?                ��/����?        ��#�� @                z�5��@                ��#�� @F�JԮDA@0#0#@��#���?��|��,@0#0#@��#���?        H�4H�4@��#���?                                H�4H�4@        ��|��,@0#0#�?        ��|��,@                        0#0#�?��#���?&jW�v%4@        ��#���?��/���@                ��/���@        ��#���?                        ��On�(@                ��/����?                �cp>'@        ��#�� @��/���@��+��+$@��#�� @��/���@H�4H�4@        ��/���@H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@        �cp>@        ��#�� @                                �C=�C=@        ��/���@�o��oyZ@        �cp>@�C=�C=@        ��/����?                ��/����?�C=�C=@                ��+��+@        ��/����?0#0# @        ��/����?                        0#0# @        0����/@_��Y��X@                �C=�C=L@        0����/@��-��-E@        �cp>@                ��/����?��-��-E@        ��/����?0#0#@        ��/����?0#0#�?                0#0#�?        ��/����?                        H�4H�4@                ��)��)C@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��NhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhMh�hhK ��h��R�(KM��h��Bh:         �                 ���?o�w�R�?3      �4� ~}@       k                  �~��?�)����?�       +�]W��u@       (                 h�"d?a����?m       �.k��d@       !                 ��??��*�K:�?&       '߫��0K@                        ��Uf?:=�����?       sl�My@@                         ��?�����?       \��j>@       
                  Pmj�?��|��?       ���ĺw@       	                 �uYJ?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               �cp>@                        @F���U�?        {|37@                        P�@?�Ug���?       ����0@                        �-�?�f%j��?       ��ꁞ9,@                        �NR?$ k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?                        h�K?p�j���?       ���z"@                        hU[U?      �<       ���>��@������������������������       �               ��#���?������������������������       �               z�5��@                        ��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?                       �-Q�f?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?                        (�&R?      �<       z�5��@������������������������       �               z�5��@������������������������       �               z�5��@                         �ȍ�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?"       #                  `���?���cE��?       c�co5@������������������������       �               ��/����?$       %                 (߁C?$#����?       w�߄�3@������������������������       �      ��       ��,���1@&       '                    �?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?)       *                 �s�?��Ԛ}�?G       n �q�[@������������������������       �               �cp>'@+       Z                 ��J?I�d���?@       &��ҩ�X@,       W                 `*�?5��>D�?/       �a��R@-       B                    �?�[�(�v�?,       |*�ӑQ@.       ;                 0�2�?�����?       r�@@/       6                  ;��?d%@�"�?       SҀh��:@0       5                 �T��?�)z� ��?       ��\�,@1       4                  �_�?x�j���?       ���z"@2       3                 ���m?����?       ��X�)B@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?������������������������       �               ;��,��@������������������������       �      ȼ       0����/@7       8                 �~�?4��c`�?       %��t5)@������������������������       �               ��/���@9       :                 (gД?, k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?<       =                  �jw?,�b���?       �GXvƒ@������������������������       �               ��#�� @>       ?                 �7��?�nɵ��?        Cad�J@������������������������       �               ��/����?@       A                 � �?�zœ���?       IG���t@������������������������       �               0#0#�?������������������������       �               z�5��@C       T                 ���?���A���?       ��\�FB@D       K                 0�?�26�
�?       6��*8E<@E       J                   .p�?xb�"���?       '�T�w1@F       G                 ���?���WW�?       �j�S@������������������������       �               z�5��@H       I                     �?���`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               \Lg1��&@L       Q                 ��e?P��W�?       94���%@M       N                   ��?r�T���?       ��e[�&@������������������������       �               ��#�� @O       P                 wu5�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?R       S                 ����?�;�a
=�?       ��l��@������������������������       �               �cp>@������������������������       �               0#0#�?U       V                 e�?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ���>��@X       Y                  �9��?<�4���?       �tCP��@������������������������       �               �cp>@������������������������       �               0#0# @[       f                 ��?v%��"�?       y=��2N8@\       ]                 ТO?��Dr�?       �9[�7�!@������������������������       �               ��/����?^       c                  �P��?���1p8�?       |곯�@_       b                  ��3�?�@����?       ���a�@`       a                 �y~?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       H�4H�4@d       e                 ���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?g       j                  ����?����VV�?	       A�R.�.@h       i                 �yQ?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �               0����/@������������������������       �               0����/#@l       �                 �2z�?_�����?x       ��P�g@m       �                    �?v�|�!�?V       �q�I+�_@n       �                  ���?���
��?:       ��V���T@o       x                 @I��>��?��?       X���F@p       q                 `���>���/��?       V��7�@������������������������       �               ��#�� @r       s                 ����?f%@�"�?       ��[�@������������������������       �               ��/����?t       u                 0?���/��?       V��7�@������������������������       �               ��#���?v       w                ppE��?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?y       ~                 @B�<?X ����?       L���B@z       {                 � }? ��vH6�?       Mߣ߶�<@������������������������       �      м       �k(��2@|       }                 NK�X?T�k����?       b*pn�$@������������������������       �               0#0#�?������������������������       �               �k(��"@       �                 �\͵?�����?       ��X�)B @������������������������       �               ��/����?������������������������       �      �<       z�5��@�       �                 0:��?���N���?       �O��!C@�       �                 @�ո?�p5Z4�?       � .J�F?@�       �                   ��?��� ��?       �{k�[=@�       �                  �E�?zp�?�r�?       �E��
$@�       �                 �o_�?�djH�E�?       ^�\m�n@�       �                 ���r?�d�$���?       �T�f@�       �                  h��?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ��#�� @�       �                   ���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               0#0#�?�       �                 ��f?Δfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@�       �                 ;��?N2o�]�?       �s��PV3@�       �                �q�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 `��~?�q���?       ��|�^1@�       �                  t�޾      �<       <��,��$@������������������������       �               ;��,��@������������������������       �               ;��,��@�       �                 ���?�)z� ��?       �\�@������������������������       �               ��#�� @�       �                 x��?
4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @������������������������       �      м       ��/����?�       �                  ?���1p8�?       |곯�@�       �                 �� �?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0#@������������������������       �               ��#���?�       �                 0)�?�Z�.�E�?       ��1�V�E@�       �                 ����?��0�Q.�?       ��c��?@�       �                 ����>x�����?       �4^$4�3@������������������������       �               ��#�� @�       �                   ��?nQ��?
       �s�=�1@������������������������       �               �cp>@�       �                 �1�?d%@�"�?       ��[�'@�       �                 �<��>      �<       ��/���@������������������������       �               ��/����?������������������������       �               �cp>@������������������������       �      ��       ��#��@�       �                 ��e|?Hj��w�?       l8�(@�       �                @5	{�?�k��?       �0QqX@������������������������       �               ��#���?������������������������       �               H�4H�4@�       �                 p�Ђ?hutee�?       Q9��@������������������������       �               0#0# @�       �                  ��d�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 �zd�?l����1�?	       ��;9�(@������������������������       �               ��#�� @������������������������       �               0#0#@�       �                 �1p�?`����r�?"       Z�c�m�L@�       �                  _��?T3��a�?       �X0�;@������������������������       �               0#0#�?�       �                 ����?jX@3��?       �(g:@�       �                 P+m�?�����f�?       4���7@������������������������       �               ���-��*@�       �                  ���?�5JH���?       �MOI#@������������������������       �               E�JԮD!@������������������������       �               0#0#�?������������������������       �               H�4H�4@�       �                 ����?S�փr�?       �+��D�=@������������������������       �               ��/����?�       �                  ���?r�7J��?       .��<@�       �                 �Q
�?(�L^{�?	       ����0&1@�       �                 ���?     ��?       "F�b@������������������������       �               H�4H�4@������������������������       �               ��#�� @�       �                  2��?v=���?       � ��R(@�       �                 �Ρ�?����|e�?       �z �B�@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?������������������������       �               0#0# @�       �                 pM�t?�it�R��?	       ��ǿ%@�       �                 �7Ө?$ k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      ��       ��/���@�       �                 `�?�?Hy��]0�?       ���y"@������������������������       �               0#0#@�       �                 ��N�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       
                 �@�?�7J�B �?N       t"M�Z�^@�                        (��?�E�+��?M       :�)�]@�       �                 h��?�(���C�?4       ��a�L6R@�       �                   �0�?���C��?#       �̕=VpH@�       �                 ��H�? �����?       C��� x-@�       �                 ����?������?       +�ǟf%@�       �                  s��?�;[��G�?       �O�;�]!@������������������������       �      �<       �cp>@�       �                 �lZ�?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �               0#0# @������������������������       �               0#0#@�       �                 �и?p��Ɵ��?       �(�NA@�       �                ���(z?      �<       �A�A>@������������������������       �        	       ��8��8*@������������������������       �               S2%S2%1@�       �                 0�2�?�@G���?       hu��@�       �                 �ޥg?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               0#0#�?�                        �6SZ?`O�+��?       j[��7@�       �                 �ڡ3?��z}-�?
       ��(�I�)@�       �                 P��?�*P��?       �����&@�       �                  `�J�?  k�Lj�?       �q��l}@������������������������       �               ��/����?�       �                 ����?`%@�"�?       ��[�@������������������������       �               ��/����?�       �                 ��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                  I��?��ڰ�x�?       �K�f�@�       �                  `s�?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?������������������������       �               z�5��@������������������������       �      ��       ��/����?                       A�?��H�&p�?       L^�3��%@������������������������       �               vb'vb'"@������������������������       �      ȼ       ��/����?                      �؉�?@`9S�?       \��Ը5G@������������������������       �               ������C@                     p�~�?�k��?       �0QqX@������������������������       �               ��+��+@      	                 =�a?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �      �       �cp>@�t�b��     h�hhK ��h��R�(KMKK��h �B  �>��d@"jW�v%d@�����b@g:��,&c@M!��a@�C=�C=L@B����R@�JԮDmS@H�4H�4(@��,���A@/����/3@        ��,���1@��/���.@        ��,���1@��On�(@        ��#�� @0����/@        ��#�� @��/����?        ��#�� @                        ��/����?                �cp>@        �P^Cy/@��/���@        �k(��"@��/���@        �k(��"@0����/@        ��#���?��/���@                ��/���@        ��#���?                ��#�� @��/����?        ���>��@                ��#���?                z�5��@                ��#���?��/����?                ��/����?        ��#���?                        �cp>@                ��/����?                ��/����?        z�5��@                z�5��@                z�5��@                        �cp>@                ��/����?                ��/����?        ��,���1@��/���@                ��/����?        ��,���1@��/����?        ��,���1@                        ��/����?                ��/����?                ��/����?        ��k(/D@H�)�BM@H�4H�4(@        �cp>'@        ��k(/D@��h
�G@H�4H�4(@������C@��|��<@�C=�C=@������C@�cp>�9@��+��+@���>��,@:l��F:2@0#0#�?�k(��"@D�JԮD1@        ��#�� @�cp>@        ��#�� @��/����?        z�5��@��/����?        z�5��@                        ��/����?        ;��,��@                        0����/@        ��#���?�cp>'@                ��/���@        ��#���?��/���@                ��/���@        ��#���?                ;��,��@��/����?0#0#�?��#�� @                z�5��@��/����?0#0#�?        ��/����?        z�5��@        0#0#�?                0#0#�?z�5��@                |�5��8@��/���@0#0#@��#��0@��/���@0#0#@���>��,@��/����?0#0# @z�5��@��/����?0#0# @z�5��@                        ��/����?0#0# @        ��/����?                        0#0# @\Lg1��&@                ��#�� @���-��@0#0# @��#�� @��/����?0#0#�?��#�� @                        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@0#0#�?        �cp>@                        0#0#�?��#�� @                ��#���?                ���>��@                        �cp>@0#0# @        �cp>@                        0#0# @��#���?:l��F:2@��+��+@��#���?��/���@0#0#@        ��/����?        ��#���?��/����?0#0#@        ��/����?0#0#@        ��/����?0#0#�?        ��/����?                        0#0#�?                H�4H�4@��#���?��/����?                ��/����?        ��#���?                        ��|��,@0#0#�?        0����/@0#0#�?                0#0#�?        0����/@                0����/#@        ���khS@2����-O@#0#0F@�k(��R@On��O@@��+��+4@    �M@D�JԮD1@�C=�C=@f:��,&C@�cp>@0#0#�?��#��@��/���@        ��#�� @                ��#�� @��/���@                ��/����?        ��#�� @��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                Ey�5A@��/����?0#0#�?+�����;@        0#0#�?�k(��2@                �k(��"@        0#0#�?                0#0#�?�k(��"@                z�5��@��/����?                ��/����?        z�5��@                <��,��4@�cp>'@H�4H�4@������3@0����/#@0#0# @������3@��/���@0#0# @;��,��@��/���@0#0#�?��#��@��/����?0#0#�?��#��@��/����?        z�5��@                ��#���?                ��#�� @                ��#���?��/����?                ��/����?        ��#���?                                0#0#�?��#���?�cp>@        ��#���?                        �cp>@        ���>��,@��/���@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?���>��,@�cp>@        <��,��$@                ;��,��@                ;��,��@                ��#��@�cp>@        ��#�� @                ��#�� @�cp>@                �cp>@        ��#�� @                        ��/����?        ��#���?��/����?0#0#@        ��/����?0#0#@        ��/����?                        0#0#@��#���?                �P^Cy/@��/���.@��8��8*@���>��@��/���.@vb'vb'"@z�5��@���-��*@        ��#�� @                ��#��@���-��*@                �cp>@        ��#��@��/���@                ��/���@                ��/����?                �cp>@        ��#��@                ��#���?��/����?vb'vb'"@��#���?        H�4H�4@��#���?                                H�4H�4@        ��/����?H�4H�4@                0#0# @        ��/����?0#0#�?                0#0#�?        ��/����?        ��#�� @        0#0#@��#�� @                                0#0#@z�5��@�_��e�=@H�4H�48@        h
��6@��+��+@                0#0#�?        h
��6@0#0#@        h
��6@0#0#�?        ���-��*@                E�JԮD!@0#0#�?        E�JԮD!@                        0#0#�?                H�4H�4@z�5��@��/���@��)��)3@        ��/����?        z�5��@�cp>@��)��)3@��#�� @��/����?�C=�C=,@��#�� @        H�4H�4@                H�4H�4@��#�� @                        ��/����?#0#0&@        ��/����?H�4H�4@                H�4H�4@        ��/����?                        0#0# @��#���?0����/@��+��+@��#���?��/���@        ��#���?                        ��/���@                ��/����?��+��+@                0#0#@        ��/����?0#0#�?        ��/����?                        0#0#�?���>��@鰑5@1��-�rW@���>��@;l��F:2@2��-�rW@z�5��@:l��F:2@H�4H�4H@        鰑%@��)��)C@        ��/���@�C=�C=@        ��/���@H�4H�4@        ��/���@0#0#�?        �cp>@                ��/����?0#0#�?        ��/����?                        0#0#�?                0#0# @                0#0#@        �cp>@=�C=�C?@                �A�A>@                ��8��8*@                S2%S2%1@        �cp>@0#0#�?        �cp>@                ��/����?                ��/����?                        0#0#�?z�5��@��/���@��+��+$@z�5��@�cp>@0#0#�?z�5��@��/���@0#0#�?��#���?��/���@                ��/����?        ��#���?��/����?                ��/����?        ��#���?��/����?                ��/����?        ��#���?                ;��,��@        0#0#�?��#�� @        0#0#�?��#�� @                                0#0#�?z�5��@                        ��/����?                ��/����?vb'vb'"@                vb'vb'"@        ��/����?        ��#���?        ;�;�F@                ������C@��#���?        H�4H�4@                ��+��+@��#���?        0#0#�?��#���?                                0#0#�?        �cp>@        �t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ2�3hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKᅔh��B81         �                 `r�t?<���G�?$      �#�,�}@       �                 `m�?b�k�9'�?�       q�A/v@                          �G�?t{��E��?�       IJcF�p@                        �R`�?R�_��?       j�͉V�H@                        p���?��Ұ��?       ��*YD@                        �,=?jy8�n�?       P(�\S'/@       
                 N���?@ǵ3���?       �q�ͨ�@       	                 ��
?r@ȱ��?       om���S@������������������������       �               0����/@������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �      ��       ��/���@                        ����?�Z�	7�?       .��9@                        @F�f����?
       $c�Z%K1@                         ��/?�3���r�?       ��7�nN*@                         ��h�j���?       ���z"@                         `s�?�����?       �O��@������������������������       �               ��/����?������������������������       �      �<       ;��,��@                        @Ws�?      �<       z�5��@������������������������       �               ��#�� @������������������������       �               ��#���?                         _4�?��fm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               ��#��@                        �Q�?̔fm���?       ��Z�N@������������������������       �      ��       �cp>@������������������������       �               ��#�� @������������������������       �               E�JԮD!@       `                 �<��?>8����?�       xS�ryk@        G                 �m�?s4M��?B       *œ�[@!       (                  �P��?�$�V��?*       ��+��Q@"       #                 @��>$#����?
       w�߄�3@������������������������       �               ��/����?$       %                 `�լ?�hK)�?	       �h��K�2@������������������������       �      ȼ       ��b:��*@&       '                 X��?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@)       B                 @B�<?l+p����?        p���XI@*       5                  ʟ�?�/�{^�?       ���B@+       0                 `���>R�䙸�?       �2	�wS7@,       -                    �?2�c3���?       �uk��!@������������������������       �               z�5��@.       /                  ;��?r@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@1       2                 ���?�DNpk�?	       �k�Z$�,@������������������������       �               z�5��(@3       4                    �?x�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?6       A                 `��?8µ*A
�?
       ��A抌)@7       @                 �饣?Ĕfm���?	       �0��z'@8       ?                 ����?���/��?       @z$S��@9       >                 eni?�Z�	7�?       j~���@:       ;                 l��w?f%@�"�?       ��[�@������������������������       �               ��/����?<       =                 @5�>���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �      м       ��/����?������������������������       �      ��       �cp>@������������������������       �      ܼ       ��#���?C       F                 p���?,0B�
��?       3j©�,-@D       E                 �<|�?h�4���?       �tCP��#@������������������������       �               �cp>@������������������������       �               0#0#@������������������������       �      ��       0����/@H       _                 pH�d?�~�Hs=�?       ,^��0rD@I       Z                 �$�?̕�z��?       .�� pC@J       Y                 �Z �?� ��i�?       �u�:hA@K       L                 P��?T�7Ke��?       �B�n�@@������������������������       �               {�5��(@M       N                 ��y�?���cE��?       c�co5@������������������������       �               ��/����?O       P                  @(B�?�3��F��?       mf9t{y4@������������������������       �               ��/����?Q       X                 ��d?$#����?       w�߄�3@R       W                 @*��?��t� �?       ����x&@S       V                 ��m?��Z�	7�?       j~���@T       U                 ����?�����?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?������������������������       �      ȼ       ��/����?������������������������       �      ��       z�5��@������������������������       �               ��#�� @������������������������       �      �<       ��/����?[       ^                 ���?|,���O�?       ���/>@\       ]                 �F��?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               0#0# @a       �                 �+@?�_!���?I       �=�@�,[@b       u                 p�%h?n��x��?*       ��#��=O@c       t                  ��ľ>hu},��?       �#�*��8@d       i                 Ш��?�Y���k�?       �b&��6@e       f                 8\Dp?�4�fP�?	       V���-@������������������������       �               ��#���?g       h                 ��V�?8��~d��?       8E���*@������������������������       �               ��On�(@������������������������       �               0#0#�?j       s                 .��U?R9�)\e�?       _���b @k       n                 (��?�_�A�?       肵�e`@l       m                  �E�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?o       r                 P�o�?�d�$���?       �T�f@p       q                 `ಣ?      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@������������������������       �      ȼ       ��/����?������������������������       �      м       ��/����?������������������������       �      �<       ��#�� @v                        ��?�N�����?       ��0�B@w       |                    �?���P��?       �*Y�ȹ9@x       {                 `�}?h�:V��?	       �GP�1@y       z                 ���?�����?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?������������������������       �               ��b:��*@}       ~                 (V�q?��6L�n�?       �E#��h @������������������������       �               ��/����?������������������������       �      �<       ���>��@�       �                 p/��?dn����?       � ��w<(@������������������������       �      м       ���>��@�       �                 �m�?  k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      �<       ��/���@�       �                 xڍ�?�J���?       �Ӟ��G@�       �                  γ�?�(Nz��?       �����E@�       �                 ��j�?p�r{��?
       e�6� /@������������������������       �               ��/���@�       �                 x8G{?Δfm���?       ��Z�N@�       �                 @� %?\n����?       � ��w<@������������������������       �               ��#���?�       �                 ��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               0����/@�       �                 ��Y?���Z�)�?       �d���;@�       �                    �?�?D] �?       #�l��8@�       �                 ��G�? ��c`�?       %��t5)@�       �                 @���?r@ȱ��?       om���S@������������������������       �               ��/���@�       �                 ��֗?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       ���-��@�       �                  ����?0�q��?	       �Mc�(@�       �                 ���?�w��d��?       �0���s@������������������������       �      �<       ��/���@������������������������       �               H�4H�4@������������������������       �      ��       ;��,��@�       �                 ��,�?      �<       z�5��@������������������������       �               ��#�� @������������������������       �               ��#���?������������������������       �      �       H�4H�4@�       �                 �{��?�ܱ�	�?:       ��:n�tU@�       �                 Ќ�j?xL�0���?       Q~�)��B@�       �                 ��a�?D_���+�?       �?�B��A@�       �                   ��?�g�vw�?       �Aws}8@������������������������       �               H�4H�4@�       �                 �j%?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?�       �                 �+#�?�g�\CY�?       A��(=@�       �                 �p�?�~���9�?       �q�Ί#6@������������������������       �      ��       ��+��+4@�       �                 ���?��G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 h6�?�Qk��?       ��Th!�@������������������������       �               �cp>@������������������������       �               0#0#@�       �                 0ɥ�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?�       �                   p��?�̥Q)�?"       <k����G@�       �                 ��Z�?
Y���a�?       �z���B@�       �                 @�t�?�A53���?       G����@@�       �                 �R�־d����?       Q	K��@�       �                  ���?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �               ��#�� @�       �                  ��?��@D�p�?       9rs~��:@�       �                    �?H�b!��?       xxZ�,�4@������������������������       �               ��#�� @�       �                 ����?��I<��?       Y���5�2@�       �                 ����?��F���?       :�.�-'@�       �                 �ſ�?$ k�Lj�?       �q��l}@������������������������       �               ��/���@������������������������       �      м       ��#���?������������������������       �               ���-��@�       �                 �ie�?�.�KQu�?       �K̎@�       �                 p���?�o���?       o�9�F@������������������������       �               ��#���?������������������������       �               0#0#@������������������������       �               ��#�� @�       �                  ���?      �<       �cp>@������������������������       �               ��/����?������������������������       �               0����/@������������������������       �               0#0#@�       �                  �{��?      �<       ��+��+$@������������������������       �               0#0#�?������������������������       �               vb'vb'"@�       �                 ��{?hm���k�?A       `qċ�c]@�       �                 n�x?p�~:��?       �����)@������������������������       �               0#0# @������������������������       �               0����/@�       �                 ��a�?��s;�?;       c2�ZK,Z@�       �                 p���?�o"����?'       ,6=i<$R@�       �                 PiU�?��4sր�?       #�	<7?@������������������������       �               �A�A>@������������������������       �      �<       ��/����?�       �                 ��=�?      �<       �ڬ�ڬD@������������������������       �               0#0#�?������������������������       �               ��+��+D@�       �                 �|_�?T�L�*��?       l���@@������������������������       �               �cp>@������������������������       �               �s?�s?=@�t�bh�hhK ��h��R�(KK�KK��h �B  y�YLGc@7l��F:b@��N�Ďe@y�YLGc@c�_��%a@Q��N��O@}�5�wa@����\@S2%S2%1@�k(��2@��/���>@        �k(��2@h
��6@        z�5��@��On�(@        z�5��@0����/@        ��#���?0����/@                0����/@        ��#���?                ��#�� @                        ��/���@        �P^Cy/@0����/#@        ��b:��*@��/���@        �k(��"@��/���@        ��#�� @��/����?        ;��,��@��/����?                ��/����?        ;��,��@                z�5��@                ��#�� @                ��#���?                ��#���?�cp>@                �cp>@        ��#���?                ��#��@                ��#�� @�cp>@                �cp>@        ��#�� @                        E�JԮD!@        r(���F^@��-��bT@S2%S2%1@j1��tVQ@�]�ڕ�?@��+��+$@d:��,&C@���-��:@��+��+@��,���1@��/����?                ��/����?        ��,���1@��/����?        ��b:��*@                ��#��@��/����?                ��/����?        ��#��@                <��,��4@��On�8@��+��+@<��,��4@��|��,@0#0#�?��#��0@�cp>@0#0#�?��#��@0����/@        z�5��@                ��#���?0����/@        ��#���?                        0����/@        z�5��(@��/����?0#0#�?z�5��(@                        ��/����?0#0#�?                0#0#�?        ��/����?        ��#��@D�JԮD!@        z�5��@D�JԮD!@        z�5��@�cp>@        z�5��@��/����?        ��#���?��/����?                ��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#�� @                        ��/����?                �cp>@        ��#���?                        鰑%@0#0#@        �cp>@0#0#@        �cp>@                        0#0#@        0����/@        �P^Cy?@0����/@��+��+@�P^Cy?@0����/@H�4H�4@Ip�}>@0����/@        Jp�}>@��/���@        {�5��(@                ��,���1@��/���@                ��/����?        ��,���1@�cp>@                ��/����?        ��,���1@��/����?        �k(��"@��/����?        z�5��@��/����?        z�5��@��/����?        z�5��@                        ��/����?                ��/����?        z�5��@                ��#�� @                        ��/����?        ��#���?        H�4H�4@��#���?        0#0#�?                0#0#�?��#���?                                0#0# @                0#0# @�#���I@��On�H@�C=�C=@��k(/D@鰑5@0#0#�?��#�� @��/���.@0#0#�?z�5��@��/���.@0#0#�?��#���?��On�(@0#0#�?��#���?                        ��On�(@0#0#�?        ��On�(@                        0#0#�?;��,��@�cp>@        ;��,��@��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#��@��/����?        ��#��@                ��#���?                z�5��@                        ��/����?                ��/����?        ��#�� @                ���b:@@�cp>@        �,����7@��/����?        ��#��0@��/����?        z�5��@��/����?        z�5��@                        ��/����?        ��b:��*@                ���>��@��/����?                ��/����?        ���>��@                ��#�� @��/���@        ���>��@                ��#���?��/���@        ��#���?                        ��/���@        [Lg1��&@��|��<@H�4H�4@[Lg1��&@��|��<@H�4H�4@��#�� @���-��*@                ��/���@        ��#�� @�cp>@        ��#�� @��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                        0����/@        �k(��"@��/���.@H�4H�4@z�5��@��/���.@H�4H�4@��#���?�cp>'@        ��#���?0����/@                ��/���@        ��#���?��/����?                ��/����?        ��#���?                        ���-��@        ;��,��@��/���@H�4H�4@        ��/���@H�4H�4@        ��/���@                        H�4H�4@;��,��@                z�5��@                ��#�� @                ��#���?                                H�4H�4@���>��,@��On�8@$S2%S2G@��#�� @��/���@�C=�C=<@��#�� @0����/@�C=�C=<@��#�� @��/����?H�4H�4@                H�4H�4@��#�� @��/����?        ��#�� @                        ��/����?                ��/���@k�6k�69@        ��/����?��-��-5@                ��+��+4@        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@0#0#@        �cp>@                        0#0#@        �cp>@                ��/����?                ��/����?        z�5��(@E�JԮD1@vb'vb'2@z�5��(@E�JԮD1@0#0# @z�5��(@D�JԮD1@0#0#@z�5��@��/����?        ��#��@��/����?        ��#��@                        ��/����?        ��#�� @                z�5��@On��O0@0#0#@z�5��@鰑%@0#0#@��#�� @                ��#��@鰑%@0#0#@��#���?鰑%@        ��#���?��/���@                ��/���@        ��#���?                        ���-��@        z�5��@        0#0#@��#���?        0#0#@��#���?                                0#0#@��#�� @                        �cp>@                ��/����?                0����/@                        0#0#@                ��+��+$@                0#0#�?                vb'vb'"@        E�JԮD!@�;�;[@        0����/@0#0# @                0#0# @        0����/@                ��/���@m�6k�6Y@        ��/����?n�fm��Q@        ��/����?�A�A>@                �A�A>@        ��/����?                        �ڬ�ڬD@                0#0#�?                ��+��+D@        �cp>@�s?�s?=@        �cp>@                        �s?�s?=@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJk�ahFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKۅ�h��B�/         �                 0V[�?	�U�B�?0      �`r}@       �                 ��y�?p�6�?��?�       �K{�kv@       �                 �6Sz?�o<ò�?�       =���r@       u                 �"��?��ʈ��?�       9nRg�p@       l                   B�?���h��?�       +����j@       C                 P�f�?��\����?       ; +Jvg@                        �$?Z?Z6[�}-�?V       �iۍ�G`@       	                 h�[�>�F���?       :�.�-7@������������������������       �               ��#���?
                        @F���/Ѷ?       ���
$6@������������������������       �        
       :l��F:2@                        @�W?Ĕfm���?       ��Z�N@                        Pkf?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��#���?       6                 ���@?XP�����?G       �(+�a�Z@       5                 ��w? V*�"�?5       iܤ?[�S@       *                 �U���Ĺ1?�V�?/       �z�Q@                        ���~?�Z�	7�?       .��9@                        ��p?�o����?	       ���5u*@                        �؉�?�����?       �O��(@������������������������       �               z�5��@                        �!�?Tn����?       � ��w<@                         <�e?`%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               z�5��@������������������������       �      м       ��/����?       '                    �?�4��v�?	       �Y-"�'@       &                 @��y?Bǵ3���?       �q�ͨ�@        !                 XΩZ?r@ȱ��?       nm���S@������������������������       �               �cp>@"       #                 ��{�?\%@�"�?       ��[�@������������������������       �               ��/����?$       %                 �dy�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#�� @(       )                 ���?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @+       ,                 � `?h����?       �Fx�v�E@������������������������       �               ��/����?-       0                 `xNv? =켴��?       �����E@.       /                  �Ԧ�?0�#�ݬ?       0X{Z�@@������������������������       �               ��/����?������������������������       �               ���b:@@1       2                 `�.8?� �_rK�?       J�@��"@������������������������       �               �cp>@3       4                  PV��?�����?       �O��@������������������������       �               ��/����?������������������������       �               ;��,��@������������������������       �               ;��,��$@7       8                 �@�?��Ұ��?       �1��<@������������������������       �               0����/#@9       >                 Ps?6�^��?       @<��*�2@:       ;                 `��z?����?       �Ä�>c(@������������������������       �               ��#�� @<       =                 ���P?Ĕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���??       @                  ��d�?�`@s'��?       Fi_y,*@������������������������       �               ��/���@A       B                 ��?h%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?D       a                  �/�?�8Ɨ}Z�?)       cEu�L@E       F                     �?�=���4�?       ��%ɡE@������������������������       �               ��/���@G       X                      &��&�?       ��Mi�A@H       O                 `��?y�!؅9�?       R���4@I       J                 �~�?��Dr�?       �9[�7�!@������������������������       �               0#0# @K       N                 0=�?l��w��?       ���@L       M                 Hq$�?$ k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?������������������������       �               0#0# @P       Q                  n:u?���Ѯ�?       ��GQ&@������������������������       �               ��/����?R       U                 0I��?h�j���?       ���z"@S       T                 ��d?      �<       ���>��@������������������������       �               ��#�� @������������������������       �               ;��,��@V       W                  ��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?Y       Z                 n�
Q?��r�S�?
       �f��%/@������������������������       �               ���-��@[       `                 ����?�`���6�?       .u��֝!@\       ]                 ��?�3`���?       .�r��@������������������������       �               0#0# @^       _                 �Eٻ?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               0����/@b       e                 �x��?�_�A�?       肵�e`,@c       d                 �3�?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@f       i                 p�T�?�FO���?	       �ߌ$@g       h                 Hq�?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ���>��@j       k                 �?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?m       r                 x�D? I��l�?       �Ȋ۫�4@n       q                 �3�_?h�:V��?
       �GP�1@o       p                 H��?\����?       P	K��@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?������������������������       �      �<       <��,��$@s       t                 �p�?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?v       �                  �~��?`=ҕ�?$       1!���(O@w       z                 `f�|?�+��*��?       �f�x*�A@x       y                 �\��?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?{       |                 ��6�?��A;�?       �����@@������������������������       �               �cp>�9@}       ~                 0Ԥ?p�r{��?       e�6� @������������������������       �               ��/���@       �                8�|�?Ɣfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?�       �                  ���?͗P����?       }t��"�:@�       �                 8���?�"6Aq�?       )$�B"@������������������������       �               ��+��+@�       �                 �e_�?�J���?       ��*]Y@������������������������       �               0#0# @������������������������       �               ��#�� @�       �                   Y��?+�� �?       gb*�}1@�       �                  P˗?,��c`�?	       %��t5)@�       �                 ��½?* k�Lj�?       �q��l}@������������������������       �               ��/����?�       �                 8��?`%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��/���@�       �                 ��2�?jutee�?       Q9��@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?�       �                 @��?�Ȯ����?       o`E\�=@������������������������       �               #0#06@�       �                  Џ~�?�Qk��?       ��Th!�@������������������������       �               H�4H�4@�       �                 X9�?�@G���?       hu��@������������������������       �               ��/����?�       �                 P�͒?z�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 0	q?�?��g��?#       �=��K�J@�       �                 @��8?��Pћ�?       M\�njm@@�       �                  v�?ڣq�t�?       ݠ/e�&3@�       �                 R|?rR����?       q\����!@�       �                 �vQ?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 ��l�?`n����?       � ��w<@������������������������       �               ��#��@������������������������       �      �<       ��/����?�       �                 @���?T,�z)(�?       H���T$@�       �                  �x��?�.�KQu�?       �K̎@������������������������       �               z�5��@������������������������       �               0#0#@������������������������       �               H�4H�4@�       �                    �?�f��!W�?       |/��&h+@�       �                 涵?�Qk��?       ��Th!�@������������������������       �               0#0#@������������������������       �               �cp>@�       �                ����?�`@s'��?       Ei_y,*@�       �                 p��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               0����/@�       �                 0��?      �<       ��+��+4@������������������������       �               H�4H�4@������������������������       �               S2%S2%1@�       �                 Ш��?����E�?I       �S0f��]@�       �                  �h?��RN���?;       l�S<W@������������������������       �               ��/����?�       �                  �g<�?(�Y���?:       �0�[p�V@�       �                    �?`H-����?       p�c#��%@�       �                 �;�?��íxq�?       $2��-�@������������������������       �               ��/���@�       �                ��D�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               ��+��+@�       �                  @���?��Z�ƽ?3       ���WQ�S@�       �                  �Mm�?��pUз?2       ��w�S@�       �                 @�-�?P�b��?"       ���"G@������������������������       �               ��8��8:@�       �                 �N��?�@����?       ���a�3@�       �                 p���?�Qk��?       ��Th!�@������������������������       �               0#0#@������������������������       �               �cp>@�       �                  �0��?�n���k�?       3��&�*@������������������������       �        	       ��+��+$@�       �                 *��?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               0#0#@@������������������������       �      �<       ��#���?�       �                 ��f?����aB�?       ��JH:@�       �                 prǥ?���ae��?	       �2��1@������������������������       �               ;��,��@�       �                 @���?)���?       T�M��)@�       �                  P���?�)z� ��?       �\�@������������������������       �               �cp>@������������������������       �               ��#��@�       �                 @w3�?�֪u�_�?       ��?�8@������������������������       �      ��       0����/@������������������������       �               0#0#�?������������������������       �               0#0# @�t�bh�hhK ��h��R�(KK�KK��h �B�  k1��tVa@�)�B�d@�fm�f�d@Ky�5�_@��z��wb@��jS@*���>�]@�]�ڕ�`@;�;�F@+���>�]@	���|�`@��)��)3@v�}w\@��]�ڕU@0#0# @�5��X@�H��tXU@H�4H�4@B����R@[�v%jWK@        ��#�� @鰑5@        ��#���?                ��#���?鰑5@                :l��F:2@        ��#���?�cp>@                �cp>@                ��/����?                ��/����?        ��#���?                ��Gp_R@�-����@@        &�}��O@��/���.@        U^CyeJ@��/���.@        �P^Cy/@/����/#@        ;��,��$@�cp>@        <��,��$@��/����?        z�5��@                ��#��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        z�5��@                        ��/����?        ;��,��@���-��@        z�5��@0����/@        ��#���?0����/@                �cp>@        ��#���?��/����?                ��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#�� @                ��#�� @��/����?                ��/����?        ��#�� @                �k(��B@�cp>@                ��/����?        �k(��B@0����/@        ���b:@@��/����?                ��/����?        ���b:@@                ;��,��@��/���@                �cp>@        ;��,��@��/����?                ��/����?        ;��,��@                ;��,��$@                ;��,��$@:l��F:2@                0����/#@        ;��,��$@E�JԮD!@        �k(��"@�cp>@        ��#�� @                ��#���?�cp>@                �cp>@        ��#���?                ��#���?�cp>@                ��/���@        ��#���?��/����?        ��#���?                        ��/����?        >��,��4@��/���>@H�4H�4@<��,��$@���-��:@H�4H�4@        ��/���@        ;��,��$@/����/3@H�4H�4@�k(��"@���-��@0#0#@��#���?��/���@0#0#@                0#0# @��#���?��/���@0#0# @��#���?��/���@                ��/���@        ��#���?                                0#0# @��#�� @�cp>@                ��/����?        ��#�� @��/����?        ���>��@                ��#�� @                ;��,��@                ��#���?��/����?                ��/����?        ��#���?                ��#���?��On�(@0#0# @        ���-��@        ��#���?�cp>@0#0# @��#���?��/����?0#0# @                0#0# @��#���?��/����?                ��/����?        ��#���?                        0����/@        <��,��$@��/���@        ��#���?�cp>@        ��#���?                        �cp>@        �k(��"@��/����?        ��#�� @                ��#���?                ���>��@                ��#���?��/����?                ��/����?        ��#���?                ��,���1@��/����?0#0# @��#��0@��/����?        z�5��@��/����?        z�5��@                        ��/����?        <��,��$@                ��#���?        0#0# @                0#0# @��#���?                ;��,��@�cp>G@#0#0&@��#�� @On��O@@0#0#�?��#���?        0#0#�?��#���?                                0#0#�?��#���?On��O@@                �cp>�9@        ��#���?���-��@                ��/���@        ��#���?�cp>@                �cp>@        ��#���?                z�5��@���-��*@��+��+$@��#�� @        �C=�C=@                ��+��+@��#�� @        0#0# @                0#0# @��#�� @                ��#���?���-��*@H�4H�4@��#���?�cp>'@        ��#���?��/���@                ��/����?        ��#���?��/����?        ��#���?                        ��/����?                ��/���@                ��/����?H�4H�4@                H�4H�4@        ��/����?                �cp>@��8��8:@                #0#06@        �cp>@0#0#@                H�4H�4@        �cp>@0#0#�?        ��/����?                ��/����?0#0#�?                0#0#�?        ��/����?        ��#�� @��On�(@0#0#@@��#�� @��On�(@H�4H�4(@���>��@��/���@0#0# @��#��@��/���@0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?        ��#��@��/����?        ��#��@                        ��/����?        z�5��@        �C=�C=@z�5��@        0#0#@z�5��@                                0#0#@                H�4H�4@��#���?D�JԮD!@0#0#@        �cp>@0#0#@                0#0#@        �cp>@        ��#���?�cp>@        ��#���?��/����?        ��#���?                        ��/����?                0����/@                        ��+��+4@                H�4H�4@                S2%S2%1@ZLg1��&@E�JԮD1@��
�pV@��#�� @/����/#@��+��+T@        ��/����?        ��#�� @��/���@��+��+T@��#���?��/���@H�4H�4@��#���?��/���@0#0#�?        ��/���@        ��#���?        0#0#�?��#���?                                0#0#�?                ��+��+@��#���?��/���@�z��z�R@        ��/���@�z��z�R@        ��/���@��-��-E@                ��8��8:@        ��/���@0#0#0@        �cp>@0#0#@                0#0#@        �cp>@                ��/����?H�4H�4(@                ��+��+$@        ��/����?0#0# @        ��/����?                        0#0# @                0#0#@@��#���?                �k(��"@��/���@vb'vb'"@�k(��"@��/���@0#0#�?;��,��@                ��#��@��/���@0#0#�?��#��@�cp>@                �cp>@        ��#��@                        0����/@0#0#�?        0����/@                        0#0#�?                0#0# @�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ6ޤhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK兔h��B2         r                 �M�?�`sPD�?,      nT�3$�}@       o                 ��?�(��z�?�       ��*<�j@       d                 �f�V?`2�r���?�       H'W��i@       !                 @Ws�?�`+�I!�?}       #Ol��gg@                        ��l�?vPc����?(       (�e}�K@                        �;�?(�Rљ�?$       ]�n��I@                         ʟ�?����?       ��w���@@                          ��?�B����?       ��<T�?@	       
                  h��?ʔfm���?       ��Z�N@������������������������       �               ��/����?                        Ǿ?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?                          ���?\�j���?       Z��\�;@                           �?�hK)�?       �h��K�2@������������������������       �      ��       ��#��0@                         �P��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?                        �5ۂ?L���'0�?       �C�� T"@������������������������       �      �<       ���>��@������������������������       �      ȼ       ��/����?                       @�~0?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��#��0@                          `���?����]L�?       N66�ͯ@                        `|)�?Ȕfm���?       ��Z�N@������������������������       �               ��/����?                       �3�.s?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               0#0#�?"       #                  ��?��ך��?U       ��&�ʆ`@������������������������       �               �cp>@$       c                 �ڡS?>���f/�?R       ŀG91�_@%       b                 ����?X�x���?P       �x��Q^@&       ?                 � �{?R�5�g�?N       �(��*�]@'       6                    �?B$�F��?'       �T��F�L@(       +                 �c�R?h�އQ�?       Շ(�fC@)       *                 �I?@ǵ3���?       �q�ͨ�@������������������������       �               0����/@������������������������       �               z�5��@,       5                  p�:?Hk� ѽ?       �����>@-       2                 G+�`?���sx�?       �iۍѧ7@.       /                 8Yt?�hK)�?       �h��K�2@������������������������       �      ��       �P^Cy/@0       1                 �j%?hn����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?3       4                 �er#?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �               ���>��@7       8                 p�V�?b!�/�'�?       t�d��"3@������������������������       �               �cp>@9       >                 �ft?X�s�	�?       e���*@:       ;                 ���r?����?       ��X�)B@������������������������       �               ��#�� @<       =                  `���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               �k(��"@@       _                 ��Ĳ?4M��1�?'       a����N@A       J                 �s�?�*f���?%       @;`��L@B       I                  �j?�}	;	�?	       uK�>4%@C       F                 P䵂?���mf�?       毠�?b@D       E                  `���?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?G       H                 ����?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               �cp>@K       P                 p��h? ��0Z��?       a��WG@L       M                    �?X�j���?       ���z"@������������������������       �               z�5��@N       O                 ��C�?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?Q       Z                 ����?:���Jx�?       �fw�M�B@R       S                 �~��?+d�^��?       ���9�J6@������������������������       �               ��|��,@T       Y                  �[�?Fǵ3���?       �q�ͨ�@U       V                 ��R�?����?       ��X�)B@������������������������       �               ��#�� @W       X                    �?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��/���@[       ^                 8�?�?^n����?	       Ԁh��K.@\       ]                 �m�?
�o����?       ���5u*@������������������������       �      ��       ;��,��$@������������������������       �      ȼ       �cp>@������������������������       �      м       ��/����?`       a                    �?      �<       ��#��@������������������������       �               z�5��@������������������������       �               ��#���?������������������������       �     ��       ��/����?������������������������       �               ;��,��@e       h                 �j�c?��4��d�?       -�V��v3@f       g                  .p�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @i       l                ����d?lO���?
       ��o0@j       k                  @��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?m       n                 ;��?��,���?       !C�s��,@������������������������       �               ���-��*@������������������������       �               0#0#�?p       q                   ҏ�?���`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0#@s       �                 @���?�l���Y�?�       �q�Fp@t       �                 ��?}
t��?u       ��ñf@u       �                 `�0z?X���O�?E       ,ݢ��Z@v       �                 �@�?���=�?5       � ͳ~T@w       �                 py?��N�?0       >6:���R@x       y                 PJ�??�Uzb,�?	       W���bn.@������������������������       �               ��+��+@z                        ����?����?       ���"�X$@{       |                 x?x�t1u�?       "�te!� @������������������������       �      ��       z�5��@}       ~                ��P}?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �      ȼ       ��/����?�       �                   ���?@�Ny�]�?'       "K8��M@�       �                 �.KR?���C�?       ��2X�B@�       �                 ��ߢ?x%��)��?       +�ڈ�>@�       �                 `U�?X ����?       2
C>�5@������������������������       �        	       ��,���1@�       �                  @mj�?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@�       �                  U��?��q�R�?       �]�{�"@�       �                 �<�?�@G���?       hu��@������������������������       �               ��/����?�       �                 �{:�?~�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                      �|2N��?       �3K}@������������������������       �               z�5��@������������������������       �               0#0# @�       �                 �!�?      �<       ���-��@������������������������       �               �cp>@������������������������       �               ��/���@�       �                 `#��?84�c�?       ]d��-�6@�       �                 p��?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?�       �                 �^�? ��k�L�?       sk��3@�       �                  � �?�L����?	       Yk���>)@�       �                 �C�J?
4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @������������������������       �               ��/���@�       �                 ���?�Qk��?       ��Th!�@�       �                 ,���?�@����?       ���a�@������������������������       �               ��/����?������������������������       �               0#0#@������������������������       �      �<       ��/����?�       �                 �߷?�;�a
=�?       ��l��@������������������������       �               0#0#�?������������������������       �               �cp>@�       �                  S)�?����9�?       �q�Ί#6@�       �                 @{ң?�?�0�!�?       a`�T�$@������������������������       �               vb'vb'"@������������������������       �      ȼ       ��/����?������������������������       �      ��	       H�4H�4(@�       �                 �N��?�D�+��?0       .N���Q@�       �                 �	I�?�ɰv��?&       Y�8�HL@�       �                 �'��?p���9��?!       � �vlH@�       �                  �9��?<V�5��?       ���u��F@������������������������       �               ��#���?�       �                   �0�?ӄ%&�?       B��>F@�       �                 p�Z?h�q����?       O�Q*s�/@�       �                  y��?�Qk��?       ��Th!�@������������������������       �               ��/����?�       �                 Ш��?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?������������������������       �               vb'vb'"@�       �                  .{�?      �<       �C=�C=<@������������������������       �               0#0#�?������������������������       �               �;�;;@�       �                 ��? �� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                    �?�~�&��?       ?�]��@������������������������       �               0#0#@�       �                 x�?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@�       �                 �81�?rqiE��?
       'aE�/@�       �                 ���?^������?       ��Iē'@�       �                 ��0�?���q���?       �:-ߩ�@�       �                   E(�?�@G���?       hu��@������������������������       �               ��/����?�       �                 x�$�?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               z�5��@������������������������       �      ��       0����/@������������������������       �               0#0#@�       �                 �xѱ?���j��?)       ��_�U@�       �                 �!�?����b�?       �{u;y�=@�       �                 P%�??�	,�?       >0�1b3@������������������������       �               �A�A.@�       �                 `��?x�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @�       �                  `���?
�
�CX�?       ��:.�%@�       �                  Z��?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#�� @������������������������       �               H�4H�4@�       �                 �;�?��e��=�?       RG-8K@�       �                 ��ݻ?8YW�m�?       ��
&(5@�       �                 ���?;�N9���?       ��{j�@�       �                 �k;�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               H�4H�4@�       �                 `B��?      �<
       0#0#0@������������������������       �               H�4H�4@������������������������       �        	       ��8��8*@������������������������       �               B�A�@@�t�bh�hhK ��h��R�(KK�KK��h �Bx  -�����d@�L!��a@׬�ڬe@��>���^@[�ڕ��T@�C=�C=@��>���^@��-��bT@H�4H�4@*���>�]@���|�P@0#0# @�k(���E@鰑%@0#0#�?���#8E@��/���@        �#���9@��/���@        �#���9@�cp>@        ��#���?�cp>@                ��/����?        ��#���?��/����?                ��/����?        ��#���?                z�5��8@�cp>@        ��,���1@��/����?        ��#��0@                ��#���?��/����?        ��#���?                        ��/����?        ���>��@��/����?        ���>��@                        ��/����?                ��/����?                ��/����?                ��/����?        ��#��0@                ��#���?�cp>@0#0#�?��#���?�cp>@                ��/����?        ��#���?��/����?                ��/����?        ��#���?                                0#0#�?C����R@�a#6�K@0#0#�?        �cp>@        B����R@��On�H@0#0#�?��,���Q@��On�H@0#0#�?��,���Q@f�_��G@0#0#�?�GpAF@���-��*@        ���b:@@���-��@        z�5��@0����/@                0����/@        z�5��@                ���>��<@��/����?        �k(���5@��/����?        ��,���1@��/����?        �P^Cy/@                ��#�� @��/����?        ��#�� @                        ��/����?        ��#��@��/����?                ��/����?        ��#��@                ���>��@                {�5��(@���-��@                �cp>@        {�5��(@��/����?        z�5��@��/����?        ��#�� @                ��#���?��/����?                ��/����?        ��#���?                �k(��"@                
�#���9@F�JԮDA@0#0#�?�k(���5@F�JԮDA@0#0#�?        /����/#@0#0#�?        ��/���@0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                �cp>@                ��/����?                ��/����?                �cp>@        �k(���5@��On�8@        ��#�� @��/����?        z�5��@                ��#�� @��/����?        ��#�� @                        ��/����?        ��b:��*@�e�_��7@        z�5��@0����/3@                ��|��,@        z�5��@0����/@        z�5��@��/����?        ��#�� @                ��#���?��/����?                ��/����?        ��#���?                        ��/���@        <��,��$@0����/@        <��,��$@�cp>@        ;��,��$@                        �cp>@                ��/����?        ��#��@                z�5��@                ��#���?                        ��/����?        ;��,��@                z�5��@��/���.@0#0#�?��#�� @��/����?                ��/����?        ��#�� @                ��#���?��|��,@0#0#�?��#���?��/����?                ��/����?        ��#���?                        ���-��*@0#0#�?        ���-��*@                        0#0#�?        ��/����?0#0#@        ��/����?                        0#0#@���#8E@R!�ML@��+��+d@������C@�e�_��G@#0#0V@��,���A@Pn��O@@xb'vb'B@��,���A@�]�ڕ�?@�A�A.@��,���A@�cp>�9@�C=�C=,@���>��@��/����?H�4H�4@                ��+��+@���>��@��/����?0#0#�?���>��@        0#0#�?z�5��@                ��#���?        0#0#�?                0#0#�?��#���?                        ��/����?        *�����;@�e�_��7@0#0# @�,����7@鰑%@H�4H�4@�,����7@��/���@H�4H�4@<��,��4@��/����?        ��,���1@                z�5��@��/����?                ��/����?        z�5��@                z�5��@�cp>@H�4H�4@        �cp>@0#0#�?        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?z�5��@        0#0# @z�5��@                                0#0# @        ���-��@                �cp>@                ��/���@        ��#��@���-��*@��+��+@��#�� @        0#0#�?��#�� @                                0#0#�?��#�� @���-��*@0#0#@��#�� @鰑%@        ��#�� @�cp>@                �cp>@        ��#�� @                        ��/���@                �cp>@0#0#@        ��/����?0#0#@        ��/����?                        0#0#@        ��/����?                �cp>@0#0#�?                0#0#�?        �cp>@                ��/����?��-��-5@        ��/����?vb'vb'"@                vb'vb'"@        ��/����?                        H�4H�4(@��#��@��/���.@��8��8J@��#���?��/���@7k�6k�G@��#���?0����/@��-��-E@��#���?�cp>@�ڬ�ڬD@��#���?                        �cp>@�ڬ�ڬD@        �cp>@��8��8*@        �cp>@0#0#@        ��/����?                ��/����?0#0#@                0#0#@        ��/����?                        vb'vb'"@                �C=�C=<@                0#0#�?                �;�;;@        ��/����?0#0#�?                0#0#�?        ��/����?                �cp>@��+��+@                0#0#@        �cp>@0#0#�?                0#0#�?        �cp>@        z�5��@��/���@��+��+@z�5��@��/���@0#0#�?z�5��@�cp>@0#0#�?        �cp>@0#0#�?        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?z�5��@                        0����/@                        0#0#@z�5��@D�JԮD!@vb'vb'R@��#�� @��/���@��+��+4@        ��/����?S2%S2%1@                �A�A.@        ��/����?0#0# @        ��/����?                        0#0# @��#�� @�cp>@H�4H�4@��#�� @�cp>@                �cp>@        ��#�� @                                H�4H�4@��#���?��/����?��8��8J@��#���?��/����?��)��)3@��#���?��/����?H�4H�4@��#���?��/����?                ��/����?        ��#���?                                H�4H�4@                0#0#0@                H�4H�4@                ��8��8*@                B�A�@@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��{hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK���h��B�)         �                 ��ݏ?�0�*T�?!      XX��؄}@       }                 ��h?��h����?�       /;�Rt@       p                   p��?f �%��?�       �ʉ2�r@       I                    �?�Gy���?�       �>�p@       
                 ��_?ӺI+���?b       �7wu��e@       	                  �^��?r@ȱ��?       ���~1@                         Z��?�h��%�?
       �1�
�u0@������������������������       �        	       ��|��,@������������������������       �               ��#�� @������������������������       �      �<       ��#���?       H                 ��?��@^�,�?W       ���C��c@       -                 @�(�?���}��?S       ��iR��b@                        ���{?(�%�K�?7       bԪ4�lZ@                        `��?PeC����?       W��_�D@                        ؝Ia?L�����?	       ��;��{5@                        ��=�?�hK)�?       �h��K�2@������������������������       �               ��,���1@������������������������       �      �<       ��/����?                        n�
Q?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?                        �>�b?      �<       �k(��2@������������������������       �               z�5��@������������������������       �        
       �P^Cy/@       $                  `��?<c�V=�?#       6����eP@                        �q�3?<St+-��?       �����E@                        �aM?jՏ�m|�?       ��h
�7@                        �o��?d%@�"�?       ��[�@������������������������       �      ��       ��/���@������������������������       �               ��#�� @������������������������       �               ��,���1@        !                 ��{�?���9��?       ����s4@������������������������       �               ���-��*@"       #                 tpx?�)z� ��?       �\�@������������������������       �               ��#��@������������������������       �               �cp>@%       (                  `s�?$c��q��?       �Y�r�5@&       '                 �aB�?��ڰ�x�?       �K�f�@������������������������       �               ;��,��@������������������������       �               0#0#�?)       *                 0I��?0k� ѽ?       �����.@������������������������       �               �k(��"@+       ,                 ���?�����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?.       C                 0i,�?䵞����?       |qP�&YF@/       B                  ���?�Z�ܙ�?       ��><QJA@0       7                  �g<�?E�$�g�?       �*XK�9@1       2                 Н@�?*I�cͿ�?	       ��J#�l'@������������������������       �               ���-��@3       4                 �lY�?��b�}�?       ���\�@������������������������       �               ��/����?5       6                 `�г?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?8       ;                 p���?{��j�?       �e��w,@9       :                 ��?�@����?       ���a�@������������������������       �               ��/����?������������������������       �               0#0#@<       ?                 @���?X�j���?       ���z"@=       >                  D&�?����?       ��X�)B@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?@       A                 ��{�?      �<       ;��,��@������������������������       �               ��#���?������������������������       �               ��#��@������������������������       �      ��       D�JԮD!@D       G                 ����?�g�(�>�?       �F�V;$@E       F                  P(B�?P�ih�<�?       ��
@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               z�5��@������������������������       �               ���-��@J       k                 8[j�?L0�[�[�?=       ?�|}�QX@K       j                  �\�?�Jz�s�?5       u$75�U@L       c                 �:W>?�_�d���?2       G�.Tk�S@M       N                 �0��>4��C��?%       ��[X)K@������������������������       �               0#0# @O       X                  �P��?������?$       ¦8('J@P       Q                  ���?&���"��?       ?8���8@������������������������       �               ��/����?R       U                 �ѱ?�ۄ���?       U:E?n�6@S       T                 @o	�? �#�Ѵ�?       �)�B�4@������������������������       �               ������3@������������������������       �      �<       ��/����?V       W                 P*�?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?Y       Z                 tlq?"$�܍�?       >R��;@������������������������       �               ��On�(@[       `                 P��?�K$e_�?       �EU�}.@\       _                 (�6�?�����?
       �O��(@]       ^                 �gZ{?ܗZ�	7�?       i~���@������������������������       �      ��       z�5��@������������������������       �      ��       ��/����?������������������������       �               ���>��@a       b                  P��?x��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @d       e                 �h!�?�L����?       Zk���>9@������������������������       �               ��/���.@f       g                 �m��?4=�%�?       �(J��#@������������������������       �               ��#�� @h       i                  ���?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#�� @������������������������       �      �       ���-��@l       o                 0\��?��H�&p�?       L^�3��%@m       n                 `ec�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0# @q       z                 ��^f?�t�Z\�?       fA�F/:@r       u                 ���?�,�_.o�?       @��*3@s       t                 Pb%�?�)z� ��?       ~�\�@������������������������       �               ��#��@������������������������       �      ȼ       �cp>@v       y                 0�H�?�/y߃�?
       ǁ\��((@w       x                  �h�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��+��+$@{       |                 0�!�?�k��?       �0QqX@������������������������       �               H�4H�4@������������������������       �               ��#���?~                        X�;�?�(�'=P�?       ( AK;@������������������������       �               ��/����?�       �                 ࢍ}?�-�bƲ?       =�7*9@������������������������       �      ��
       vb'vb'2@�       �                 X�)�?d�ih�<�?       ��
@������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?�       �                 �$�c?+l����?]       ��S�db@�       �                 �' �?����p��?&       a�n �O@�       �                 p�-�?�d�$���?       �T�f$@������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?�       �                 �d|�?���*��?!       -��u��J@�       �                 0�C�?�J���?       ���t�o$@�       �                 PJ�?��ڰ�x�?       �K�f�@������������������������       �               ;��,��@������������������������       �               0#0#�?������������������������       �               0#0#@�       �                 ��*�?�Ei��?       m�X��E@�       �                 �Ψ?�֪u�_�?       ��?�8'@������������������������       �               ���-��@�       �                 ����?`�4���?       �tCP��@������������������������       �               �cp>@������������������������       �               0#0# @�       �                   �0�?T��0�z�?       ����?@�       �                 ����?>b����?       �}IS6@�       �                 ��?Ȕfm���?       ��Z�N@������������������������       �               ��#�� @������������������������       �               �cp>@�       �                  p%+�?~��j�?	       �e��w,@������������������������       �               ��/����?�       �                 `�>?T����1�?       ��;9�(@�       �                  ��?��$4��?       �F�.Tk"@�       �                 pMH�?��h��?       S�D'�@������������������������       �               ��#��@�       �                 ���?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               0#0# @������������������������       �      ȼ       z�5��@�       �                 PeT�?����h�?       @��o{#@������������������������       �               0#0# @�       �                  p��?xLU���?       i�ҹ^�@�       �                 ���H?      �<       ���-��@������������������������       �               ��/���@������������������������       �               �cp>@������������������������       �               0#0#�?�       �                  ��d�? ���h�?7       �o6�T@�       �                    �?.�4��?       p��P9�0@������������������������       �               H�4H�4@�       �                 ���?��Ñp��?       <7��0�%@�       �                  @��?|��`p��?       f;3@��!@������������������������       �               0#0#@�       �                 Pl?l�4���?       �tCP��@������������������������       �               0#0#�?�       �                 ��B�?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �      м       ��/����?�       �                 p�:�?�~���9�?,       `����P@�       �                  ~�?�j.�d��?       �I���+@�       �                    �?x�G���?       '5L�`�@������������������������       �               H�4H�4@������������������������       �               �cp>@������������������������       �               0#0# @������������������������       �      ��!       ��8��8J@�t�b��     h�hhK ��h��R�(KK�KK��h �B�  ��k(/d@/����/c@������c@YUUUU5a@u�����]@M�dJ��P@YUUUU5a@=�)�B]@�
��
�E@�,���n`@L!�M\@�;�;;@�5��X@Qn��OP@��8��8*@z�5��@��|��,@        ��#�� @��|��,@                ��|��,@        ��#�� @                ��#���?                ����JW@n��F:lI@��8��8*@����JW@h
��F@��8��8*@�b:���S@�e�_��7@0#0# @�YLg1B@�cp>@0#0#�?��,���1@�cp>@0#0#�?��,���1@��/����?        ��,���1@                        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?�k(��2@                z�5��@                �P^Cy/@                �k(���E@鰑5@0#0#�?�,����7@%jW�v%4@        ������3@��/���@        ��#�� @��/���@                ��/���@        ��#�� @                ��,���1@                ��#��@On��O0@                ���-��*@        ��#��@�cp>@        ��#��@                        �cp>@        ������3@��/����?0#0#�?;��,��@        0#0#�?;��,��@                                0#0#�?���>��,@��/����?        �k(��"@                ;��,��@��/����?        ;��,��@                        ��/����?        ��b:��*@'jW�v%4@#0#0&@;��,��$@0����/3@��+��+@<��,��$@鰑%@��+��+@��#�� @D�JԮD!@0#0#�?        ���-��@        ��#�� @��/����?0#0#�?        ��/����?        ��#�� @        0#0#�?��#�� @                                0#0#�?��#�� @��/����?0#0#@        ��/����?0#0#@        ��/����?                        0#0#@��#�� @��/����?        z�5��@��/����?        z�5��@                        ��/����?        ;��,��@                ��#���?                ��#��@                        D�JԮD!@        z�5��@��/����?H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@z�5��@                        ���-��@        ��,���A@�e�_��G@�C=�C=,@��,���A@�cp>G@��+��+@��,���A@������C@��+��+@�P^Cy?@;l��F:2@��+��+@                0#0# @�P^Cy?@:l��F:2@H�4H�4@;��,��4@�cp>@0#0#�?        ��/����?        ;��,��4@��/����?0#0#�?������3@��/����?        ������3@                        ��/����?        ��#���?        0#0#�?                0#0#�?��#���?                <��,��$@��/���.@0#0# @        ��On�(@        <��,��$@�cp>@0#0# @<��,��$@��/����?        z�5��@��/����?        z�5��@                        ��/����?        ���>��@                        ��/����?0#0# @        ��/����?                        0#0# @��#��@鰑5@                ��/���.@        ��#��@�cp>@        ��#�� @                ��#�� @�cp>@                �cp>@        ��#�� @                        ���-��@                ��/����?vb'vb'"@        ��/����?0#0#�?                0#0#�?        ��/����?                        0#0# @z�5��@��/���@0#0#0@;��,��@��/���@��+��+$@��#��@�cp>@        ��#��@                        �cp>@        ��#���?��/����?��+��+$@��#���?��/����?                ��/����?        ��#���?                                ��+��+$@��#���?        H�4H�4@                H�4H�4@��#���?                        �cp>@H�4H�48@        ��/����?                ��/����?H�4H�48@                vb'vb'2@        ��/����?H�4H�4@                H�4H�4@        ��/����?        �,����7@�-����@@��
�pV@�,����7@�cp>�9@�C=�C=,@��#�� @��/����?        ��#�� @                        ��/����?        �P^Cy/@�e�_��7@�C=�C=,@;��,��@        ��+��+@;��,��@        0#0#�?;��,��@                                0#0#�?                0#0#@<��,��$@�e�_��7@vb'vb'"@        0����/#@0#0# @        ���-��@                �cp>@0#0# @        �cp>@                        0#0# @<��,��$@��|��,@�C=�C=@;��,��$@��/���@0#0#@��#�� @�cp>@        ��#�� @                        �cp>@        ��#�� @��/����?0#0#@        ��/����?        ��#�� @        0#0#@;��,��@        0#0#@;��,��@        0#0# @��#��@                ��#���?        0#0# @��#���?                                0#0# @                0#0# @z�5��@                        ���-��@H�4H�4@                0#0# @        ���-��@0#0#�?        ���-��@                ��/���@                �cp>@                        0#0#�?        ��/���@�i��R@        0����/@H�4H�4(@                H�4H�4@        0����/@H�4H�4@        �cp>@H�4H�4@                0#0#@        �cp>@0#0# @                0#0#�?        �cp>@0#0#�?        �cp>@                        0#0#�?        ��/����?                �cp>@P��N��O@        �cp>@#0#0&@        �cp>@H�4H�4@                H�4H�4@        �cp>@                        0#0# @                ��8��8J@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ?{�hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKυ�h��BH-         l                 @@�?��W�4�?*      ���Kz}@       c                  �a�?bf+X��?�       �k�#�k@       P                 0��?� �1��?�       όu��i@       E                 ���@?���o���?h       �'�:e@       "                 )DW?DZ��M��?T       Ç��a@                        @��l?^�A ��?/       ��7e�;R@                        ���L?�4��v�?       �Y-"�7@������������������������       �               ��#��@	                        @F�~�����?       �4^$4�3@
                        `�t$?�(�����?       ��0��0@                        �aH�>|���A�?       /gX\-@������������������������       �               ��#�� @������������������������       �        	       ��On�(@                       @`�e&?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?                        `%�7?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?       !                 pt"?(FX}Q2�?       �7³��H@                        8Yt?��b�J��?       ��?��>@                        `��?X ����?       2
C>�5@                        �k�J?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@                        ,*���      �<       ��#��0@������������������������       �               ��#�� @������������������������       �               ���>��,@                        ��Ɲ?j%@�"�?       �6�E�!@������������������������       �               �cp>@                            �?      �<       z�5��@������������������������       �               ��#�� @������������������������       �               ��#���?������������������������       �        
       �k(��2@#       .                 P^s?��pp?+�?%       {�שIQ@$       %                 ��-�?��\���?       �̑-`R9@������������������������       �               ��#�� @&       -                    �?t�r{��?       �)i@7@'       (                 ���>f%@�"�?       �6�E�!@������������������������       �               �cp>@)       ,                 M}?���/��?       @z$S��@*       +                 XJ��?�Z�	7�?       j~���@������������������������       �               z�5��@������������������������       �      �<       ��/����?������������������������       �      м       ��/����?������������������������       �      ��       ��|��,@/       B                 �Y�b?�����?       y�<�E@0       7                  �v�?u�����?       ��r�K@@1       2                  �"�?�	�����?
       Yr��9�3@������������������������       �               z�5��@3       4                 @�6{?إ�je��?	       ��BLGh0@������������������������       �      �<       ��On�(@5       6                  ��?z�G���?       ��%�|@������������������������       �               0#0# @������������������������       �      �<       ��/����?8       ?                 �T�?@�d��N�?	       =��g�%*@9       :                 �>œ?bn����?       ~��Y-"@������������������������       �      ��       ;��,��@;       <                 �(�?Ȕfm���?       ��Z�N@������������������������       �               ��#���?=       >                 �ܝ�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?@       A                  Pmj�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@C       D                 �/��?��t� �?       ����x&@������������������������       �               �k(��"@������������������������       �      ȼ       ��/����?F       I                  `��?�ZKގ��?       ';d�:@G       H                 0�?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?J       O                 �Z�?�B�� �?       �HI�7@K       L                  ���?�F���?	       :�.�-'@������������������������       �      ��       ��/���@M       N                 ���?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �      �<	       �cp>'@Q       Z                 �ڬ�?F8�e�?       H��}UMB@R       W                 �R�־��6L�n�?       ��4}i�8@S       V                    �?<9�)\e�?       _���b @T       U                 ��?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               ��#��@X       Y                ��W�y?      �<
       ��#��0@������������������������       �               ��b:��*@������������������������       �               z�5��@[       b                 ��(�?�\U�?	       �{����'@\       a                 ��|?���`�?       ��
�Me@]       ^                  �"�?l@ȱ��?       om���S@������������������������       �      �<       ��/���@_       `                 ����?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               ��#��@d       i                 ��;�?B������?
       ��6�س0@e       f                 G҈n?�'z�3�?       ���da�%@������������������������       �               ��+��+@g       h                 ����?�� ��?       qp� k@������������������������       �               0#0# @������������������������       �      ��       ��/���@j       k                 tՀ�?�֪u�_�?       ��?�8@������������������������       �               0����/@������������������������       �               0#0#�?m       �                 ����?-PK�!/�?�       ��r�Fo@n       �                 @��`?�fs���?x       Q;ɼ5\g@o       �                    �? x$�?D       Rn^�*�X@p       q                   ���?z�,����?'       D��@�M@������������������������       �               D�JԮD!@r       �                 ��N�?>哧I��?"       �%�-�I@s       t                 x��?�>Q0�8�?       ���g��F@������������������������       �               H�4H�4@u       ~                  ����?X�N����?       T�z3XzE@v       {                 P&��?�w͘�?       �I����*@w       x                 �Um�?d7Y���?	       ���r�&@������������������������       �               �k(��"@y       z                  ���?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?|       }                 ��i�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?       �                 ����?v���ߡ�?       г"�=@�       �                 3^�?���y���?       D��$�9@�       �                  `���?��"��b�?
       _���d�2@������������������������       �               0����/@�       �                 ��f�?�.4�v��?       &�~F�,@������������������������       �               z�5��@�       �                  ��?V����?       �Y9��%@������������������������       �               ��/����?�       �                 �i�?��q�R�?       �]�{�"@�       �                 �C�J?b,���O�?       ���/>@������������������������       �               H�4H�4@������������������������       �               ��#���?�       �                  0���?
4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @�       �                  p��?<�a
=�?       ��l��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �               0#0#@�       �                 P��?      �<       ;��,��@������������������������       �               ��#���?������������������������       �               ��#��@�       �                 @��?зH5��?       e��C@������������������������       �               ��/���@�       �                 0'�[?k;�$��?       ���H�@@�       �                 ��?�χ�O�?       )����'?@�       �                  �a�?��6L�n�?       �E#��h @������������������������       �               ��#��@�       �                 'uk?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@�       �                 ����?v���;)�?       B��"Z�6@�       �                  �.�?X�ih�<�?       W�3D*5@������������������������       �               ��/����?�       �                �I�s?�?�0�!�?       a`�T�4@������������������������       �      ��       #0#0&@�       �                  �9��?h����?       �����!@������������������������       �               0#0# @�       �                 0?�AP�9��?       h��6��@������������������������       �               ��/����?������������������������       �      ��       ��+��+@�       �                 ��x�?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �      �<       ��/����?�       �                 ��9�?dɮ����?4       T4�@�U@�       �                 ��c�?������?3       �H��tXU@�       �                 @2i�?�ƛO�?+       �e�aR@�       �                  M}�?8f��{�?       ��C&=@������������������������       �               0#0#0@�       �                 �y�?�N�+�?
       ����*@�       �                  �a�?v=���?	       � ��R(@������������������������       �               ��/����?������������������������       �               #0#0&@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       #0#0F@�       �                 ��?��ό��?       ���C��'@������������������������       �               ��/����?�       �                 �^��?*^�yU�?       ��7�1�#@������������������������       �               ��+��+@�       �                 ��j�?l�4���?       �tCP��@�       �                 �5��?z��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �      �<       ��/����?������������������������       �      �<       ��/����?�       �                 �؉�?����?&       n��T�O@�       �                   E(�?�ɮ����?#       r`E\�M@������������������������       �               �cp>@�       �                 0�Ь?ع�f
@�?!       "?uG�K@�       �                 P%�?����|e�?       7\@��'@�       �                p��ש?�?�0�!�?       a`�T�$@�       �                 P��?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0# @������������������������       �      ȼ       ��/����?������������������������       �      ��       �
��
�E@�       �                  �2�?��|2N��?       �3K}@������������������������       �               z�5��@������������������������       �               0#0# @�t�bh�hhK ��h��R�(KK�KK��h �Bh  YUUUU5a@鰑Nc@
��
�pf@V^CyeZ@�D�J�.Y@�A�A.@V^CyeZ@�cp>W@�C=�C=@������S@鰑U@��+��+@f:��,&S@;��18N@��+��+@V^CyeJ@&jW�v%4@        <��,��$@���-��*@        ��#��@                z�5��@���-��*@        ��#��@��On�(@        ��#�� @��On�(@        ��#�� @                        ��On�(@        ��#�� @                ��#���?                ��#���?                ��#�� @��/����?        ��#�� @                        ��/����?        ���#8E@���-��@        �,����7@���-��@        <��,��4@��/����?        ��#��@��/����?                ��/����?        ��#��@                ��#��0@                ��#�� @                ���>��,@                z�5��@�cp>@                �cp>@        z�5��@                ��#�� @                ��#���?                �k(��2@                �,����7@'jW�v%D@��+��+@;��,��@%jW�v%4@        ��#�� @                z�5��@%jW�v%4@        z�5��@�cp>@                �cp>@        z�5��@�cp>@        z�5��@��/����?        z�5��@                        ��/����?                ��/����?                ��|��,@        �k(��2@&jW�v%4@��+��+@�k(��"@:l��F:2@��+��+@z�5��@��|��,@0#0# @z�5��@                        ��|��,@0#0# @        ��On�(@                ��/����?0#0# @                0#0# @        ��/����?        z�5��@��/���@H�4H�4@z�5��@�cp>@        ;��,��@                ��#���?�cp>@        ��#���?                        �cp>@                ��/����?                ��/����?                ��/����?H�4H�4@        ��/����?                        H�4H�4@�k(��"@��/����?        �k(��"@                        ��/����?        ��#�� @�e�_��7@        ��#���?��/����?                ��/����?        ��#���?                ��#���?h
��6@        ��#���?鰑%@                ��/���@        ��#���?�cp>@                �cp>@        ��#���?                        �cp>'@        ��b:��:@��/���@0#0# @�k(���5@�cp>@        ;��,��@�cp>@        ��#���?�cp>@                �cp>@        ��#���?                ��#��@                ��#��0@                ��b:��*@                z�5��@                ;��,��@0����/@0#0# @��#���?0����/@0#0# @��#���?0����/@                ��/���@        ��#���?��/����?                ��/����?        ��#���?                                0#0# @��#��@                        E�JԮD!@0#0# @        ��/���@�C=�C=@                ��+��+@        ��/���@0#0# @                0#0# @        ��/���@                0����/@0#0#�?        0����/@                        0#0#�?���b:@@���-��J@ȔLɔ�d@���>��<@�e�_��G@�����{[@���>��<@������C@=�C=�C?@�k(���5@��On�8@��8��8*@        D�JԮD!@        �k(���5@On��O0@��8��8*@��#��0@On��O0@��8��8*@                H�4H�4@��#��0@On��O0@��+��+$@<��,��$@��/����?0#0# @<��,��$@        0#0#�?�k(��"@                ��#���?        0#0#�?                0#0#�?��#���?                        ��/����?0#0#�?        ��/����?                        0#0#�?z�5��@��/���.@0#0# @z�5��@��/���.@0#0#@z�5��@0����/#@H�4H�4@        0����/@        z�5��@0����/@H�4H�4@z�5��@                z�5��@0����/@H�4H�4@        ��/����?        z�5��@�cp>@H�4H�4@��#���?        H�4H�4@                H�4H�4@��#���?                ��#�� @�cp>@                �cp>@        ��#�� @                        �cp>@0#0#�?        �cp>@                        0#0#�?                0#0#@;��,��@                ��#���?                ��#��@                ���>��@��|��,@vb'vb'2@        ��/���@        ���>��@���-��@vb'vb'2@���>��@�cp>@vb'vb'2@���>��@��/����?        ��#��@                z�5��@��/����?                ��/����?        z�5��@                        0����/@vb'vb'2@        �cp>@vb'vb'2@        ��/����?                ��/����?vb'vb'2@                #0#0&@        ��/����?�C=�C=@                0#0# @        ��/����?��+��+@        ��/����?                        ��+��+@        ��/����?                ��/����?                ��/����?                ��/����?                E�JԮD!@������S@        ���-��@������S@        ��/����?n�fm��Q@        ��/����?�;�;;@                0#0#0@        ��/����?#0#0&@        ��/����?#0#0&@        ��/����?                        #0#0&@        ��/����?                        #0#0F@        0����/@�C=�C=@        ��/����?                �cp>@�C=�C=@                ��+��+@        �cp>@0#0# @        ��/����?0#0# @                0#0# @        ��/����?                ��/����?                ��/����?        z�5��@�cp>@�;�;K@        �cp>@��8��8J@        �cp>@                �cp>@��8��8J@        �cp>@vb'vb'"@        ��/����?vb'vb'"@        ��/����?0#0#�?                0#0#�?        ��/����?                        0#0# @        ��/����?                        �
��
�E@z�5��@        0#0# @z�5��@                                0#0# @�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��}whFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK酔h��B�2         �                 p��?>��:+M�?,      �Յi	}@       �                  t0�?��:�?      ��vu�{@       �                 �8U|?�ul#�?�       �L�[xu@       q                   �x�?B���%��?�       ���jes@       Z                  �~��?�q&���?�       �u�"��i@       ;                 �c=d?�,��.�?^       X[��a@       .                  �P��?P=���J�?=       l�_�V@                        ��f?��1���?1       �� [��R@	                        (+�g?Z�'��?       ��2�D@
                        �U����#�1o�?       hI"炵?@                        X��?<9�)\e�?       _���b @������������������������       �               �cp>@������������������������       �               ;��,��@                        @��>��sx�?       �iۍѧ7@������������������������       �               ��/����?                        ���}?�(1k��?       �ꁞ9�6@������������������������       �               \Lg1��&@                        ��c�?����X��?       &��֞&@������������������������       �               ��/����?������������������������       �               ;��,��$@                        J�e?���/��?       5��o��#@������������������������       �               ;��,��@������������������������       �      ��       0����/@       +                  �9��?x�$/^%�?       �_���@@       *                   .p�?�R�u-��?       .=kD\=@                        �a ?Par[+Z�?       i!�Y<@������������������������       �               ��#���?                        �m�?xf�T6|�?       {,*��P;@������������������������       �               �cp>'@                        Z�K?Bǵ3���?       �q�ͨ�/@������������������������       �               ��#���?        #                 p���?`%@�"�?       ̰rɱ�-@!       "                ��U%�?��Z�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@$       )                 P�s�?& k�Lj�?       �q��l}#@%       &                 �b��?b%@�"�?       ��[�@������������������������       �               ��#���?'       (                 ����?$ k�Lj�?       �q��l}@������������������������       �      �<       ��/���@������������������������       �               ��#���?������������������������       �      ��       ��/���@������������������������       �               0#0#�?,       -                 0�3%?      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@/       :                 ���P?��fm���?       ��Z�N/@0       5                   s��?&µ*A
�?	       ��A抌)@1       2                 (�?�`@s'��?       Fi_y,*@������������������������       �               ��#���?3       4                 `s5�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               0����/@6       7                 �yW?���/��?       @z$S��@������������������������       �               ��/����?8       9                    �?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@������������������������       �               �cp>@<       W                 0�2�?����zP�?!       L2��I@=       F                   ��?�:��$�?       t�6�E�G@>       ?                 �Q�?� ����?       �	��+9@������������������������       �      ��	       鰑5@@       C                 ��=�?����?       ��X�)B@A       B                 xT2P?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?D       E                    �?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?G       L                 Pώ?IU����?       "��N��5@H       K                 ���m?���Ѯ�?       ��GQ&@I       J                 8�4b?���/��?       @z$S��@������������������������       �               �cp>@������������������������       �               z�5��@������������������������       �      �<       ;��,��@M       T                      ^�ђ���?
       �oFݜh%@N       O                    �?
4=�%�?       �(J��@������������������������       �               ��#���?P       Q                  @?��?Ȕfm���?       ��Z�N@������������������������       �               ��#���?R       S                  p�~?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?U       V                 `u?      �<       �cp>@������������������������       �               ��/����?������������������������       �               0����/@X       Y                  �G?�?      �<       z�5��@������������������������       �               ��#�� @������������������������       �               ��#���?[       d                 ���@?�zV�w�?%       ;#O�P@\       c                 p^��?�G|:=*�?       �`���G@]       b                  ���?J)�$fz�?       �Ulz�x9@^       _                 Б{�?�fB��?
       �^q�,,@������������������������       �               ��#�� @`       a                 0��?�֪u�_�?       ��?�8@������������������������       �               0����/@������������������������       �               0#0#�?������������������������       �               ZLg1��&@������������������������       �        
       �k(���5@e       n                 ��o�?�� :��?       �*�b��2@f       m                  ��d�?���/��?       J9U6�+@g       l                    �?0k�"O��?       �?<��*&@h       k                  ~��?jP�D�?       �A��P?$@i       j                  �Q�?F���'0�?       �C�� T"@������������������������       �               ��/����?������������������������       �               ���>��@������������������������       �      м       ��/����?������������������������       �      м       ��/����?������������������������       �      Լ       �cp>@o       p                 `�.�?hutee�?       Q9��@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?r       �                 p'v�?*+��Tc�?;       #��*�Y@s       �                 `��?!�!4�?4       ��I�J2V@t       �                 `�Hj?�&��ռ�?       ��~���?@u       �                 �]t?ĸ�qA��?       �����5@v       }                    �?�d�$���?
       <��#�.@w       x                 �$y=?|b8�Y�?       EJͰ(@������������������������       �               ���>��@y       |                 _�
?~d�$���?       �T�f@z       {                 p��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      �<       z�5��@~                        ��/?b%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                  �:D?�֪u�_�?       ��?�8@������������������������       �               0����/@������������������������       �               0#0#�?�       �                 �.��?�^�#΀�?       O�{��A%@������������������������       �               0����/#@������������������������       �      ܼ       ��#���?�       �                 ����?T�p�@/�?        ��S�L@�       �                 �p�?��X����?       ⳱���E@�       �                 @5�>�pe�(p�?       ����D@�       �                  pjS�?z��`p��?       ��u��4@�       �                 ��?l�K�+:�?       �ޖ��2@�       �                  ��^�?��Ñp��?       <7��0�%@������������������������       �               �cp>@�       �                ��z?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               0#0# @������������������������       �      м       ��/����?�       �                  �G?�?w�%
�j�?       JQlČ-3@�       �                 ���?)�ť��?       Z`Il�7,@������������������������       �               ���>��@�       �                    �?�w��d��?       �0���s@������������������������       �               �cp>@�       �                 @���?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                P3��`?�o���?       o�9�F@�       �                   ���?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               H�4H�4@�       �                 ����?      �<       ��/���@������������������������       �               ��/����?������������������������       �               �cp>@�       �                 p/��?�S��W��?	       $$�
�g*@������������������������       �               �k(��"@�       �                  `s�?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@�       �                 Hoۆ?��&���?       ��G2��,@�       �                ���ms?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��On�(@�       �                    �?H�N�u�?       i���@@������������������������       �      ��       S2%S2%1@�       �                  �E�?w�;B��?
       ՟���	0@�       �                  LG�?�AP�9��?       h��6��@�       �                 ��;�?Hy��]0�?       ���y"@������������������������       �               ��+��+@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?������������������������       �               vb'vb'"@�       �                  �g<�?t��� �?D       /�bi�X@�       �                 Ш��?�^���?       ?P��9@�       �                 ��?�'z�3�?       ���da�%@�       �                 ��?�� ��?       rp� k@������������������������       �               0#0# @������������������������       �      �<       ��/���@������������������������       �               ��+��+@�       �                 �1ݧ?�_�A�?       炵�e`,@�       �                 ��=�?�����?       �O��(@������������������������       �      �<       <��,��$@������������������������       �      ȼ       ��/����?������������������������       �      м       ��/����?�       �                 p�f�?�����?5       ����R@�       �                  P�"�?D��NV=�?       �t�ܲ@������������������������       �               ��/����?�       �                    �?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?�       �                   p��? u��?2       �	�Y�Q@�       �                 `�4x?��`c���?&       �v�J@�       �                 p=�?��ʜ#�?       fy���6@������������������������       �               0#0#@�       �                  �Ԧ�?�n�]:��?       ٸ����2@�       �                 `�>?�D#���?       �B�j@������������������������       �               0#0#@������������������������       �               ��#�� @�       �                 ���? @�����?	       \n\�/V)@������������������������       �               ��/���@�       �                 0C�?�����?       �v�qp�!@�       �                  �^��?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?������������������������       �      ��       ��/���@������������������������       �               �s?�s?=@������������������������       �               vb'vb'2@�       �                 ��|�? [���G�?       � `0?)=@�       �                 ؗ�j?��r��?       D?J�]3@�       �                 �s�?�*P��?       �����&@�       �                  ���?���A���?       ��\�F"@������������������������       �               ��#��@�       �                 ���?��b�}�?       ���\�@�       �                 �t_�?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?�       �                  `���?w�;B��?       ՟���	 @������������������������       �               H�4H�4@�       �                 8��?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��+��+$@�t�bh�hhK ��h��R�(KK�KK��h �B�  -�����d@�B�)Dd@wb'vb'b@�����c@������c@V��N��_@�YLg1b@ 6�aca@	����M@�YLg1b@e�_��%a@�C=�C=<@Sg1��4\@���|NV@��+��+@���b:P@t�'�x�R@0#0#�?�,����G@鰑E@0#0#�?�k(���E@��/���>@0#0#�?���b:@@0����/#@        ��b:��:@0����/@        ;��,��@�cp>@                �cp>@        ;��,��@                �k(���5@��/����?                ��/����?        �k(���5@��/����?        \Lg1��&@                ;��,��$@��/����?                ��/����?        ;��,��$@                ;��,��@0����/@        ;��,��@                        0����/@        \Lg1��&@鰑5@0#0#�?���>��@鰑5@0#0#�?���>��@鰑5@        ��#���?                z�5��@鰑5@                �cp>'@        z�5��@0����/#@        ��#���?                ;��,��@/����/#@        z�5��@��/����?                ��/����?        z�5��@                ��#�� @��/���@        ��#�� @��/���@        ��#���?                ��#���?��/���@                ��/���@        ��#���?                        ��/���@                        0#0#�?��#��@                ��#���?                z�5��@                ��#��@�cp>'@        ��#��@D�JԮD!@        ��#���?�cp>@        ��#���?                        �cp>@                ��/����?                0����/@        z�5��@�cp>@                ��/����?        z�5��@��/����?                ��/����?        z�5��@                        �cp>@        ��#��0@�-����@@        ��b:��*@�-����@@        z�5��@h
��6@                鰑5@        z�5��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                ��#���?                ��#���?                <��,��$@�cp>'@        ��#�� @�cp>@        z�5��@�cp>@                �cp>@        z�5��@                ;��,��@                ��#�� @D�JԮD!@        ��#�� @�cp>@        ��#���?                ��#���?�cp>@        ��#���?                        �cp>@                ��/����?                ��/����?                �cp>@                ��/����?                0����/@        z�5��@                ��#�� @                ��#���?                6��tSH@���-��*@0#0#@>��,��D@0����/@0#0#�?������3@0����/@0#0#�?��#�� @0����/@0#0#�?��#�� @                        0����/@0#0#�?        0����/@                        0#0#�?ZLg1��&@                �k(���5@                ���>��@E�JԮD!@H�4H�4@���>��@���-��@        ���>��@��/���@        ���>��@�cp>@        ���>��@��/����?                ��/����?        ���>��@                        ��/����?                ��/����?                �cp>@                ��/����?H�4H�4@                H�4H�4@        ��/����?        ���b:@@�e�_��G@%S2%S27@�P^Cy?@E�JԮDA@%S2%S27@��b:��*@D�JԮD1@0#0#�?{�5��(@��/���@0#0#�?z�5��(@�cp>@        [Lg1��&@��/����?        ���>��@                ��#��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        z�5��@                ��#���?��/����?        ��#���?                        ��/����?                0����/@0#0#�?        0����/@                        0#0#�?��#���?0����/#@                0����/#@        ��#���?                ��,���1@D�JԮD1@#0#06@��#�� @��|��,@��-��-5@��#�� @鰑%@��-��-5@        ���-��@�C=�C=,@        0����/@�C=�C=,@        0����/@H�4H�4@        �cp>@                ��/����?H�4H�4@        ��/����?                        H�4H�4@                0#0# @        ��/����?        ��#�� @��/���@�C=�C=@���>��@��/���@H�4H�4@���>��@                        ��/���@H�4H�4@        �cp>@                ��/����?H�4H�4@        ��/����?                        H�4H�4@��#���?        0#0#@��#���?        0#0#�?                0#0#�?��#���?                                H�4H�4@        ��/���@                ��/����?                �cp>@        �k(��"@�cp>@0#0#�?�k(��"@                        �cp>@0#0#�?                0#0#�?        �cp>@        ��#���?���-��*@        ��#���?��/����?                ��/����?        ��#���?                        ��On�(@                ��/����?=�C=�C?@                S2%S2%1@        ��/����?�C=�C=,@        ��/����?��+��+@        ��/����?��+��+@                ��+��+@        ��/����?                ��/����?                        vb'vb'"@��b:��*@:l��F:2@L�dJ��P@;��,��$@��/���@�C=�C=@        ��/���@�C=�C=@        ��/���@0#0# @                0#0# @        ��/���@                        ��+��+@<��,��$@��/���@        ;��,��$@��/����?        <��,��$@                        ��/����?                ��/����?        z�5��@鰑%@�A�AN@��#���?��/����?0#0#�?        ��/����?        ��#���?        0#0#�?��#���?                                0#0#�?��#�� @D�JԮD!@����M@��#�� @E�JԮD!@�ڬ�ڬD@��#�� @D�JԮD!@H�4H�4(@                0#0#@��#�� @E�JԮD!@0#0# @��#�� @        0#0#@                0#0#@��#�� @                        E�JԮD!@0#0#@        ��/���@                0����/@0#0#@        ��/����?0#0#@                0#0#@        ��/����?                ��/���@                        �s?�s?=@                vb'vb'2@z�5��@0����/@vb'vb'2@z�5��@0����/@0#0# @z�5��@��/���@0#0#�?z�5��@��/����?0#0#�?��#��@                ��#�� @��/����?0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?��#�� @                        ��/����?                ��/����?�C=�C=@                H�4H�4@        ��/����?0#0#�?        ��/����?                        0#0#�?                ��+��+$@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�,�hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKӅ�h��B(.         �                  /Ⱥ?V��BHH�?(      �D�Ή}@       a                 ���?Ь��d3�?�       �ǐ�f�p@       H                 0G?�ot��-�?�       ������j@       ;                 0>~?�_�G��?o       t,J��e@                        �\ͥ?̔*�0 �?Z       ��j�`@                        � �5?�C=+��?       b��T|0@������������������������       �               ��/����?������������������������       �      ��       �P^Cy/@	       
                  ���?ܬ�Q%��?N       �ۅ��H]@������������������������       �               ���>��@       ,                 ����?��cos�?L       �җ�y[@       !                 ,*���̕9�/�?8       w�.;S@                         �u��?2��u��?       ��4}�A@������������������������       �               ���-��@                        �ìW?:�����?       �^��=@                         �"�?N�ђ���?       �oFݜh%@������������������������       �               ��/���@                         x�>��|��?       ���ĺw@������������������������       �               ��#���?                        hH�??r@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@                         p5W�?�����?       N��o�g2@                        ���g?�x�<�?       X&b��q1@������������������������       �               ��#�� @                         Џ~�?B���'0�?       �C�� T"@������������������������       �      �<       ;��,��@                        P��?���/��?       V��7�@������������������������       �               ��/����?                         `s�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      �<       ��/����?"       +                   ��?�FO���?       	�ߌD@#       $                 �5�?�����?       ��X�)B0@������������������������       �               ��#�� @%       (                  @(B�?���/��?       V��7�@&       '                 xux?�����?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?)       *                 $�4?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �      ��       |�5��8@-       0                  �9��?�p���K�?       E2(ߪ{@@.       /                 ��?h�4���?       �tCP��@������������������������       �               0#0# @������������������������       �               �cp>@1       :                 h�B?nw��?       c�?�-<@2       5                  L��?��F��^�?       Ҧ (2	;@3       4                  ;��?h�4���?       �tCP��@������������������������       �               �cp>@������������������������       �               0#0# @6       9                 �]��>��/Ѷ?       ���
$6@7       8                 ��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �        
       %jW�v%4@������������������������       �      �<       ��#���?<       A                  �9��?��+��?       ���|��C@=       @                    �?�)z� ��?       �\�@>       ?                 ��O1?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               z�5��@B       C                 ��N�?�C=+��?       c��T|@@������������������������       �               ������3@D       G                 �If�?�(߫$��?       1H����*@E       F                 8���?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               �k(��"@I       Z                  `%+�?\c�`�N�?       ���K�D@J       S                   s��?�?8�խ�?       ��A�7>@K       P                 ��F�?�}>D�P�?       �狢G5@L       O                 ��I?������?       �N0gX1@M       N                 P<�\?& k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      �<       ��/���@������������������������       �      �<       ��On�(@Q       R                 ��`m?|�G���?       ��%�|@������������������������       �               0#0# @������������������������       �      �<       ��/����?T       Y                  ~��?8�c3���?       �uk��!@U       X                 `��?^n����?       � ��w<@V       W                 T��?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �               �cp>@[       `                 n�
Q?Ң��'�?       �^��$@\       ]                 8} Q?f%@�"�?       ��[�@������������������������       �               ��/����?^       _                 ��l?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               �C=�C=@b       s                    �?��[���?'       ����a�L@c       p                 ����?�s ��?       -$�H�=@d       o                  f?� ����?       �趩��3@e       j                 ��f�?���6�?       0Oi]q)@f       g                 0N��?��b�}�?       ���\�@������������������������       �               ��/����?h       i                 ����?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?k       n                 �_�?hLU���?       i�ҹ^�@l       m                 ཥ�?      �<       ���-��@������������������������       �               �cp>@������������������������       �               ��/���@������������������������       �               0#0#�?������������������������       �               �C=�C=@q       r                  `<��?�?�0�!�?       a`�T�$@������������������������       �               vb'vb'"@������������������������       �      ȼ       ��/����?t       w                 �༡? &4�X �?       �(�z�;@u       v                 �s�?�����?       �O��@������������������������       �      �<       ;��,��@������������������������       �      ȼ       ��/����?x                        P:;�?��R�z�?        Gwr��5@y       ~                 0vb�?n-�E�T�?       ��<)@z       }                 `ݭ�?����|e�?       �z �B�@{       |                 �&��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               0#0# @������������������������       �      ��       E�JԮD!@�       �                 �ߦx?�iE���?        ��_�8"@�       �                  E(�?�_�A�?       肵�e`@������������������������       �               ��/����?������������������������       �               ;��,��@������������������������       �               0#0# @�       �                 �4�?���qR�?u       ����"i@�       �                 ����?��\0�?6       ���T@�       �                 p��{?��צ��?       ��,[ufE@�       �                  �9��?����w�?       L�A5ٴ?@������������������������       �               E�JԮD!@�       �                    �?�|V<���?       �]ˁ7@�       �                  �Ԡ?,Lj����?       ���T�@������������������������       �               z�5��@������������������������       �               0#0#�?�       �                 ��n�?����w�?       G�A5ٴ/@�       �                 @xA�?�*P��?       �����&@������������������������       �               ��#��@�       �                 ��{?�Z�ܙ�?       d����@������������������������       �               ��/���@�       �                 �@��?X����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �      ȼ       0����/@������������������������       �               #0#0&@�       �                 �N��?����
�?       4�r�^D@�       �                   �0�?�}+�Ҽ�?       [�B5"�8@�       �                  Ц6�?h�4���?       �tCP��#@�       �                 ~R�?z��`p��?       �����@�       �                 �~�?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �               H�4H�4@������������������������       �      �<       ��/���@������������������������       �      �<
       �A�A.@�       �                 ��j�?vqiE��?
       'aE�/@������������������������       �               0����/@�       �                 0am�?+�oI���?       ~�V&@�       �                   ��?Ȕfm���?       ��Z�N@������������������������       �               ��#���?�       �                 ���?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?�       �                  Џ~�?��3Fi�?       :�"Ξs@������������������������       �               ��#�� @������������������������       �               ��+��+@�       �                 �Nͼ?N��д�??       ���>�b]@�       �                 ���?����e�?       ���3@@�       �                ����?��P����?       <#��,@ @�       �                 �j%?����|e�?       �z �B�@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?������������������������       �               ��#��@�       �                  ���?\,���0�?       �гkQ8@�       �                 p�L�?`���X��?	       Oà4�42@������������������������       �               �A�A.@�       �                ����?H����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?�       �                 �!�?~�G���?       '5L�`�@������������������������       �               H�4H�4@������������������������       �               �cp>@�       �                 �xѱ?��=�
�?-       ^�K�SU@�       �                 �!�?�!���?       Yt<k{@@�       �                 p�/c?D�b��?	       ���"7@������������������������       �               H�4H�4(@�       �                 �)�?��H�&p�?       L^�3��%@�       �                ��ǎ�?lutee�?       Q9��@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �      ��       H�4H�4@�       �                 ��V�?熛���?       �7vg�#@������������������������       �               ��/���@�       �                 _%?��]ۀ��?       E���O@�       �                 �*�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               0#0#@�       �                  ~�?��s;�?       b2�ZK,J@�       �                 0Dh�?����|e�?       �z �B�@������������������������       �               ��+��+@�       �                  \��?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �      ��       #0#0F@�t�bh�hhK ��h��R�(KK�KK��h �B�  ��b:��c@Z<�œb@�~��~ne@�5�װ`@h��F:lY@vb'vb'B@s(���F^@h
���S@��8��8*@��P^C�\@Z�v%jWK@0#0#@�b:���S@��On�H@0#0#@�P^Cy/@��/����?                ��/����?        �P^Cy/@                ���b:P@z%jW�vH@0#0#@���>��@                w�}wL@x%jW�vH@0#0#@�>��nK@h
��6@        ��,���1@:l��F:2@                ���-��@        ��,���1@�cp>'@        ��#�� @E�JԮD!@                ��/���@        ��#�� @0����/@        ��#���?                ��#���?0����/@        ��#���?                        0����/@        �P^Cy/@�cp>@        �P^Cy/@��/����?        ��#�� @                ���>��@��/����?        ;��,��@                ��#�� @��/����?                ��/����?        ��#�� @��/����?                ��/����?        ��#�� @                        ��/����?        �k(��B@��/���@        |�5��(@��/���@        ��#�� @                ��#��@��/���@        z�5��@��/����?        z�5��@                        ��/����?        ��#���?�cp>@                �cp>@        ��#���?                |�5��8@                ��#�� @���-��:@0#0#@        �cp>@0#0# @                0#0# @        �cp>@        ��#�� @�e�_��7@0#0# @��#���?�e�_��7@0#0# @        �cp>@0#0# @        �cp>@                        0#0# @��#���?鰑5@        ��#���?��/����?        ��#���?                        ��/����?                %jW�v%4@        ��#���?                ��,���A@0����/@        ��#��@�cp>@        ��#���?�cp>@                �cp>@        ��#���?                z�5��@                �P^Cy?@��/����?        ������3@                [Lg1��&@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        �k(��"@                z�5��@��On�8@vb'vb'"@;��,��@�cp>7@0#0# @��#���?9l��F:2@0#0# @��#���?On��O0@        ��#���?��/���@        ��#���?                        ��/���@                ��On�(@                ��/����?0#0# @                0#0# @        ��/����?        ��#��@0����/@        ��#��@��/����?        ��#��@��/����?                ��/����?        ��#��@                        ��/����?                �cp>@        ��#���?��/����?�C=�C=@��#���?��/����?                ��/����?        ��#���?��/����?        ��#���?                        ��/����?                        �C=�C=@z�5��(@h
��6@%S2%S27@��#�� @/����/#@vb'vb'2@��#�� @E�JԮD!@vb'vb'"@��#�� @E�JԮD!@0#0# @��#�� @��/����?0#0#�?        ��/����?        ��#�� @        0#0#�?��#�� @                                0#0#�?        ���-��@0#0#�?        ���-��@                �cp>@                ��/���@                        0#0#�?                �C=�C=@        ��/����?vb'vb'"@                vb'vb'"@        ��/����?        <��,��$@��On�(@��+��+@;��,��@��/����?        ;��,��@                        ��/����?        ;��,��@�cp>'@��+��+@        0����/#@H�4H�4@        ��/����?H�4H�4@        ��/����?0#0#�?        ��/����?                        0#0#�?                0#0# @        E�JԮD!@        ;��,��@��/����?0#0# @;��,��@��/����?                ��/����?        ;��,��@                                0#0# @[Lg1��6@��]�ڕE@K�dJ��`@�P^Cy/@��/���>@�z��z�B@z�5��(@E�JԮD1@��8��8*@{�5��(@E�JԮD1@0#0# @        E�JԮD!@        {�5��(@E�JԮD!@0#0# @z�5��@        0#0#�?z�5��@                                0#0#�?z�5��@D�JԮD!@0#0#�?z�5��@��/���@0#0#�?��#��@                ��#�� @��/���@0#0#�?        ��/���@        ��#�� @        0#0#�?                0#0#�?��#�� @                        0����/@                        #0#0&@z�5��@���-��*@H�4H�48@        �cp>@��)��)3@        �cp>@0#0#@        ��/����?0#0#@        ��/����?0#0#�?        ��/����?                        0#0#�?                H�4H�4@        ��/���@                        �A�A.@z�5��@��/���@��+��+@        0����/@        z�5��@�cp>@��+��+@��#���?�cp>@        ��#���?                        �cp>@                ��/����?                ��/����?        ��#�� @        ��+��+@��#�� @                                ��+��+@���>��@��On�(@T�PuX@z�5��@��/���@#0#06@��#��@��/����?H�4H�4@        ��/����?H�4H�4@                H�4H�4@        ��/����?        ��#��@                ��#�� @�cp>@��)��)3@��#�� @        0#0#0@                �A�A.@��#�� @        0#0#�?��#�� @                                0#0#�?        �cp>@H�4H�4@                H�4H�4@        �cp>@        ��#���?D�JԮD!@�i��R@��#���?���-��@k�6k�69@        ��/����?��-��-5@                H�4H�4(@        ��/����?vb'vb'"@        ��/����?H�4H�4@        ��/����?                        H�4H�4@                H�4H�4@��#���?0����/@0#0#@        ��/���@        ��#���?��/����?0#0#@��#���?��/����?                ��/����?        ��#���?                                0#0#@        ��/����?n�6k�6I@        ��/����?H�4H�4@                ��+��+@        ��/����?0#0#�?                0#0#�?        ��/����?                        #0#0F@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�%\hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKم�h��Bx/         �                  ɉ�?��Ek=P�?(      �v5�e�}@       �                 0�0�?@n���?�       ���a��t@       h                 �.��?��.���?�       @j�D:q@       U                 ��?2p��D/�?z       ���ä�g@       B                 ���@?��)z���?b       �Ȑ�?c@       3                 �U����N���?L       jLd�$`@       $                    �?��xS+�?1       �̓>��S@                        �"R?����?        ��J�xJ@	       
                  �a�?��Xv#�?       )RҀh�4@������������������������       �               E�JԮD!@                        p���>�4��v�?       �Y-"�'@������������������������       �               z�5��@                        �/��?nQ��?       �s�=�!@                       ��r?l�r{��?       e�6� @������������������������       �               ���-��@������������������������       �               ��#���?������������������������       �               ��#���?                         L��?&7*��=�?       �Õ��?@                         ��g�?0�(��?       ��V-�:@������������������������       �               ��/����?                        �I?̝�/U��?       �+�f��9@                        ���?H�'e��?       �F�ҽn0@������������������������       �      ��       \Lg1��&@                        P��s?ҟ��X�?       l�n�/@                        p�^�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?                        �~�?R����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �               �k(��"@        !                  �P�? k�Lj�?       �q��l}@������������������������       �               ��/����?"       #                 ���?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?%       0                   ��?B�왓�?       �^y��g:@&       /                 P�^�?A
:����?       {��"�%@'       (                 �7�<?���/��?       5��o��#@������������������������       �               �cp>@)       .                  h��?�_�A�?       肵�e`@*       -                 ���`?�����?       �O��@+       ,                   .p�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ��       z�5��@������������������������       �      ȼ       ��/����?������������������������       �               0#0#�?1       2                 �Ux�?�Tu��?	       ����.@������������������������       �               ��|��,@������������������������       �      �<       ��#���?4       ?                 �:W>?��٤���?       � �H@5       >                 ����?����>?�?       �vD���F@6       7                 PhaX?����?       F����F@������������������������       �               0����/@8       ;                 ���p? �$3�i�?       ��7���C@9       :                 �r?��=�Sο?       ����,@������������������������       �               ��b:��*@������������������������       �      ȼ       ��/����?<       =                 pŔ�>      �<       |�5��8@������������������������       �               z�5��@������������������������       �               �k(���5@������������������������       �      �<       ��/����?@       A                 �#�?4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @C       R                   ���?S�@�~�?       ��cq9@D       O                 �6��?f��M�?       7B��	�2@E       J                 Pc	�?>ĩAf�?       ��d>v�0@F       G                 @F�e��}�?       ��Se+@������������������������       �        
       鰑%@H       I                 h��?^%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?K       L                 0A��?��q�R�?       C}Ԥ@������������������������       �               ��#���?M       N                 ׻�s?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?P       Q                 �M�s?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?S       T                 �W�V?d�ih�<�?       ��
@������������������������       �               ��/����?������������������������       �               H�4H�4@V       W                 0��}?��o�J��?       ��A8B@������������������������       �               ��|��,@X       _                 0vb�?�a�ێ
�?       �n�|W6@Y       ^                 @vn�?�)w�q�?       ��|��-@Z       [                 �5W�?v=���?	       � ��R(@������������������������       �               �C=�C=@\       ]                 @rk?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       �cp>@`       a                  χ�?���j�?       �e��w@������������������������       �               0#0#�?b       c                 �N<�?�djH�E�?       ^�\m�n@������������������������       �               z�5��@d       e                 ��P�?��q�R�?       C}Ԥ@������������������������       �               ��#���?f       g                 P}�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?i       j                 ��D?(��Z��?1       ⟆���T@������������������������       �               0����/@k       �                 n�?�2�D�g�?0       .�V��vS@l       �                 ����?�n�9��?#       ����M@m       �                 `}��?�>A��?"       ��T�x�L@n       u                 ��\�?�!:de�?        +�&ޔ�K@o       r                  ���?��?	       ��l}�'*@p       q                 
kol?j��H��?       v�I�@������������������������       �               z�5��@������������������������       �      ��       ��/���@s       t                 �m�?�����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?v       w                 �[1)?=켴��?       �����E@������������������������       �               ��/����?x       �                 ��{�?�FO���?       �ߌD@y       ~                 ����?�@US�?       �g�l�9@z       }                   �G�?X ����?       0
C>�5@{       |                ��W�y?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��	       ������3@       �                �3�q?̔fm���?       ��Z�N@������������������������       �               ��/����?�       �                 `U�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               �P^Cy/@�       �                    �?j�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 �se?��"��b�?       `���d�2@�       �                 �'+�?��z}-�?       ��(�I�)@�       �                 �jU?C�pB}��?       ����1$@�       �                 �\��?$Lj����?       ���T�@������������������������       �               ;��,��@�       �                 p%�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �      ȼ       �cp>@�       �                 PFe�?�� ��?       qp� k@�       �                 �5Ry?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      ��       �cp>@�       �                 p۶�?=���E�?'       k)��LN@�       �                 �$�c?�DHf�?       6@��zA@�       �                 ���?��íxq�?	       $2��-�'@�       �                 ��´?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @�       �                 ��0�?�(���?       y��uk!@�       �                 ��W�?f%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �      �<       �cp>@�       �                 �\ͥ?      �<       %S2%S27@������������������������       �               0#0# @������������������������       �               ��-��-5@�       �                 ��p?x(MbȎ�?       �i��g�9@������������������������       �               ��/����?�       �                 Dm�p?�zœ���?       ��x�Ϯ8@������������������������       �               �k(��2@������������������������       �               H�4H�4@�       �                 ����?
�����?V       Ѿ�"Ma@�       �                 ��l`?R96�Q�?Q       ��z(�5`@�       �                 @Y��?H��)���?'       H�;�LL@�       �                 ���H?.I�ML�?       ia���?@�       �                  ���?�rh�.��?       ����6@�       �                   �x�?�%E�N��?       �h���2@�       �                 ����?���_`�?       &!j�\+"@�       �                 ��0�?ܗZ�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@�       �                  �a�?b,���O�?       ���/>@������������������������       �               ��#���?������������������������       �               H�4H�4@�       �                 0���?���mf�?       寠�?b#@�       �                  `���?�;[��G�?       �O�;�]!@�       �                    �?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ���-��@������������������������       �               0#0#�?������������������������       �               ��#��@�       �                    �?      �<       E�JԮD!@������������������������       �               �cp>@������������������������       �               �cp>@�       �                 `�(�?��W���?       "���9@�       �                 �6SZ?�w��d��?       �0���s@������������������������       �      �<       ��/���@������������������������       �               H�4H�4@�       �                  0�?��^�}�?       �d�-.2@������������������������       �               ��#���?������������������������       �               S2%S2%1@�       �                    �?��Yk���?*       C��KER@������������������������       �               �;�;;@�       �                 PiU�?-��ޭ�?       ��	�F@������������������������       �               ��+��+$@�       �                  ��?��%O���?       ��Z�A@������������������������       �               ��/���@�       �                 0�=�?�́[B�?       #,����?@�       �                  �x��?t}��e��?       Z���0@������������������������       �               ��+��+@�       �                 p}c�?�!�a6Z�?       ���t0�'@������������������������       �               ��+��+@������������������������       �               ���-��@������������������������       �        	       �A�A.@�       �                �g�?���^���?       ���w!@������������������������       �               0#0# @������������������������       �      ��       ���-��@�t�b�t     h�hhK ��h��R�(KK�KK��h �BX  ,�����d@g
���c@�4H�4�b@���khc@v�����]@�s?�s?M@#�}��`@�a#6�[@�;�;;@>��,��T@鰑U@%S2%S27@������S@Rn��OP@��+��+$@B����R@��On�H@H�4H�4@��,���A@&jW�v%D@H�4H�4@���>��<@鰑5@0#0# @;��,��@��/���.@                E�JԮD!@        ;��,��@���-��@        z�5��@                ��#�� @���-��@        ��#���?���-��@                ���-��@        ��#���?                ��#���?                �,����7@�cp>@0#0# @\Lg1��6@��/����?0#0# @        ��/����?        \Lg1��6@��/����?0#0# @��b:��*@��/����?0#0# @\Lg1��&@                ��#�� @��/����?0#0# @        ��/����?0#0#�?        ��/����?                        0#0#�?��#�� @        0#0#�?                0#0#�?��#�� @                �k(��"@                ��#���?��/���@                ��/����?        ��#���?��/����?        ��#���?                        ��/����?        z�5��@/����/3@0#0#�?;��,��@0����/@0#0#�?;��,��@0����/@                �cp>@        ;��,��@��/����?        ;��,��@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                z�5��@                        ��/����?                        0#0#�?��#���?��|��,@                ��|��,@        ��#���?                ��k(/D@/����/#@        e:��,&C@���-��@        f:��,&C@�cp>@                0����/@        e:��,&C@��/����?        ��b:��*@��/����?        ��b:��*@                        ��/����?        |�5��8@                z�5��@                �k(���5@                        ��/����?        ��#�� @�cp>@                �cp>@        ��#�� @                z�5��@��/���.@�C=�C=@z�5��@��|��,@0#0#�?��#�� @���-��*@0#0#�?��#���?��On�(@                鰑%@        ��#���?��/����?                ��/����?        ��#���?                ��#���?��/����?0#0#�?��#���?                        ��/����?0#0#�?                0#0#�?        ��/����?        ��#���?��/����?        ��#���?                        ��/����?                ��/����?H�4H�4@        ��/����?                        H�4H�4@��#��@0����/3@��8��8*@        ��|��,@        ��#��@0����/@��8��8*@        ��/���@#0#0&@        ��/����?#0#0&@                �C=�C=@        ��/����?0#0#@                0#0#@        ��/����?                �cp>@        ��#��@��/����?0#0# @                0#0#�?��#��@��/����?0#0#�?z�5��@                ��#���?��/����?0#0#�?��#���?                        ��/����?0#0#�?                0#0#�?        ��/����?        �#���I@���-��:@0#0#@        0����/@        �#���I@h
��6@0#0#@\Lg1��F@��On�(@0#0#�?^Lg1��F@鰑%@0#0#�?\Lg1��F@0����/#@        ��#�� @0����/@        z�5��@��/���@        z�5��@                        ��/���@        ;��,��@��/����?        ;��,��@                        ��/����?        �k(��B@0����/@                ��/����?        �k(��B@��/���@        �k(���5@��/���@        <��,��4@��/����?        ��#���?��/����?                ��/����?        ��#���?                ������3@                ��#���?�cp>@                ��/����?        ��#���?��/����?        ��#���?                        ��/����?        �P^Cy/@                        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?        z�5��@/����/#@H�4H�4@z�5��@�cp>@0#0#�?z�5��@�cp>@0#0#�?z�5��@        0#0#�?;��,��@                ��#���?        0#0#�?��#���?                                0#0#�?        �cp>@                �cp>@                ��/���@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @        �cp>@        <��,��4@D�JԮD!@=�C=�C?@��#�� @��/���@k�6k�69@��#�� @��/���@0#0# @��#���?        0#0# @��#���?                                0#0# @��#���?��/���@        ��#���?��/����?                ��/����?        ��#���?                        �cp>@                        %S2%S27@                0#0# @                ��-��-5@�k(��2@��/����?H�4H�4@        ��/����?        �k(��2@        H�4H�4@�k(��2@                                H�4H�4@�k(��"@������C@��
�pV@�k(��"@On��O@@��o���U@�k(��"@h
��6@k�6k�69@��#�� @:l��F:2@��+��+@��#�� @0����/#@��+��+@��#��@/����/#@��+��+@��#��@��/����?H�4H�4@z�5��@��/����?                ��/����?        z�5��@                ��#���?        H�4H�4@��#���?                                H�4H�4@        ��/���@0#0# @        ��/���@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        ���-��@                        0#0#�?��#��@                        E�JԮD!@                �cp>@                �cp>@        ��#���?��/���@��+��+4@        ��/���@H�4H�4@        ��/���@                        H�4H�4@��#���?        S2%S2%1@��#���?                                S2%S2%1@        鰑%@>�C=�CO@                �;�;;@        鰑%@dJ�dJ�A@                ��+��+$@        鰑%@k�6k�69@        ��/���@                ���-��@k�6k�69@        ���-��@��+��+$@                ��+��+@        ���-��@��+��+@                ��+��+@        ���-��@                        �A�A.@        ���-��@0#0# @                0#0# @        ���-��@        �t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ2�hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKÅ�h��B�*         �                 ��g? �TC�=�?&      w?d��}@       y                 (�?�'�[Ę�?�       �d!9�v@       ^                 �� <?(�ݬ�?�       ]df�p@       Q                 ����?�'Y�=�?w       ���c��j@       P                 0>~?�DV�h��?j       ����Rg@       E                  �v�?"���Hr�?\       �J�"�d@       @                 �xK�?���7�T�?J       ��N�%_@       +                    �?Z��=��?A       FH��~[@	                        �U����L�]�?+       �A�E#~R@
                        �3}?�O�y���?       }����A@                          ��?��x�5��?       ���|�@@������������������������       �               �cp>@                        ���m?��h!��?       X�v%jW;@                        pae?����ɚ�?       �^��!5@                        ��?������?       +x�1�)@                        `��?�Z�	7�?       j~���$@                        0�Q�?f%@�"�?       ��[�@                        �؉�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ��       �cp>@������������������������       �               ��#��@������������������������       �      Լ       �cp>@                        p��h?��6L�n�?       �E#��h @������������������������       �      �<       ���>��@������������������������       �      ȼ       ��/����?                        0�?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ;��,��@������������������������       �      �       �cp>@       (                 �8�?L���m>�?       1w��e�B@        %                 x��?��0��5�?       �8���A@!       "                 `�]?`�s�	�?       e���*@������������������������       �               ��#�� @#       $                 ��?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?&       '                 �Z��>      �<       �k(���5@������������������������       �               ��#���?������������������������       �               <��,��4@)       *                  ��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?,       7                 ��p?���ae��?       �2��A@-       4                 ��� ?��/ʪ��?       G�Ų��1@.       1                  Џ~�?� �_rK�?       J�@��"@/       0                 �;�?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@2       3                �>�o.?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@5       6                 .25Q?      �<       D�JԮD!@������������������������       �               �cp>@������������������������       �               �cp>@8       ;                 ���5?�G�.>�?       tDB��Y2@9       :                 ��{?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@<       =                 h�?0Lj����?       ���T�,@������������������������       �               <��,��$@>       ?                 ���?�J���?       ��*]Y@������������������������       �               0#0# @������������������������       �               ��#�� @A       D                  �T? k�Lj�?	       e*�}#<-@B       C                  >�?l��H��?       v�I�@������������������������       �               ��/���@������������������������       �      �<       z�5��@������������������������       �      �<       ��/���@F       M                 �T�?�^O<.��?       �P;�B@G       L                 ��`�?��+�*�?       wȚ�
A@H       K                 �2�:?\����?       P	K��@I       J                 �j%?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               ��#��@������������������������       �      ��       ��b:��:@N       O                 �b�?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               �#���9@R       S                  +�?H�Q-���?       ��P�n;@������������������������       �               0#0#@T       U                 `�?3y�d��?       ^�1f7@������������������������       �               ��#���?V       Y                 ;��?��a���?
       �>�A6]6@W       X                   E(�?lutee�?       Q9��@������������������������       �               ��/����?������������������������       �               H�4H�4@Z       [                 @��?)���?       y��uk1@������������������������       �               E�JԮD!@\       ]                 ��s'?jQ��?       �s�=�!@������������������������       �               ���-��@������������������������       �               ��#�� @_       r                 кI�?�=EƢ��?#       �7���uI@`       a                 `�b?Z�ђ���?       �oFݜhE@������������������������       �               0����/#@b       o                 @�ޅ?�(�����?       ��0��@@c       d                 ��vi?����A�?       2gX\=@������������������������       �               ��#�� @e       f                 P��?e��}�?       ��Se;@������������������������       �        
       ��On�(@g       h                  t:t?t���A�?
       0gX\-@������������������������       �               ��#���?i       l                  ���?e��}�?	       ��Se+@j       k                 ����?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?m       n                  |1q?      �<       0����/#@������������������������       �               ��/����?������������������������       �               ��/���@p       q                  ����?      �<       ��#��@������������������������       �               ��#�� @������������������������       �               ��#�� @s       t                 Б4�?z��x���?       �!��4 @������������������������       �               ��#��@u       x                 �^7�?D��NV=�?       �t�ܲ@v       w                 (vb�?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �      �<       ��/����?z       �                   p��?����2P�?B       �-�J�CX@{       �                 pOA�?4��G�?2       �Tk��S@|       �                 Ш��?��Ml��?#       Ċ&���K@}       �                 �fů?h�4���?       �tCP��3@~       �                 `ec�?r�~:��?       �����)@       �                 @E��?���};��?
       ��;̑�%@�       �                 �jE?h�4���?       �tCP��@������������������������       �               0#0# @������������������������       �               �cp>@������������������������       �      ��       H�4H�4@������������������������       �      м       ��/����?������������������������       �      ��       ���-��@�       �                  �Q�?�l@5�q�?       r��t)B@������������������������       �               ;��,��$@�       �                 A��?�O����?       F۔m�9@�       �                 �3��?H�b!��?       xxZ�,�4@�       �                 `/D�?�F�?!�?       2V���2@������������������������       �               0#0# @�       �                 �@�?��߭Q��?
       �QVl�0@�       �                 0�C�?R�ђ���?       �oFݜh%@������������������������       �      ��       E�JԮD!@������������������������       �               ��#�� @�       �                  `���?\n����?       � ��w<@������������������������       �               ��#��@������������������������       �      �<       ��/����?������������������������       �               0#0# @������������������������       �      ؼ       ;��,��@�       �                  ���?N��Σ4�?       >`�� 7@�       �                  �X�?�˷���?       ���4��#@�       �                   �P�?�ǧ\�?       �,W J@������������������������       �               0����/@������������������������       �               H�4H�4@������������������������       �               ��#�� @������������������������       �               ��8��8*@�       �                  �{��?      �<       vb'vb'2@������������������������       �               H�4H�4@������������������������       �               �A�A.@�       �                  ��~�?(����<�?J       SKx���[@������������������������       �               ��#�� @�       �                 `��?��nd��?I       �X�>I[@������������������������       �               ��/����?�       �                    �?$�l]��?H       ���r�Z@������������������������       �               ��+��+D@�       �                 �2��?>)>:Ċ�?*       ,:����P@�       �                 ���?���fņ�?       ҋ�'8@�       �                 ާ�?d*�'=P�?        �2"@�       �                  ����?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               ��+��+@������������������������       �      ��	       �A�A.@�       �                 ���?��N�t�?       J��-]E@�       �                 P���? �Ϟi�?       ��RE�:@�       �                 �4��?*^�yU�?       ��7�1�3@�       �                 ����?h�4���?       �tCP��@������������������������       �               ��/����?�       �                  9ר?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                  ����?�@����?
       	}M��-@������������������������       �               0#0# @�       �                 0~?�Qk��?       ��Th!�@������������������������       �               ��/����?�       �                 �Ր�?�@����?       ���a�@�       �                  �0��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       H�4H�4@�       �                 \�ϸ?<�a
=�?       ��l��@������������������������       �               �cp>@������������������������       �               0#0#�?�       �                 ��e�?`r����?	       Qz�i0@������������������������       �      ��       �A�A.@������������������������       �      ȼ       ��/����?�t�bh�hhK ��h��R�(KK�KK��h �BH  �GpAf@z����a@�i��b@�#����e@��`@�[��[�L@U^Cyc@k��F:lY@#0#0&@k1��tVa@Pn��OP@��+��+$@5��t�`@�e�_��G@H�4H�4@�>��n[@ f�_��G@H�4H�4@B����R@��h
�G@0#0# @�YLg1R@����z�A@0#0# @��b:��J@&jW�v%4@        ������3@Nn��O0@        ������3@���-��*@                �cp>@        ������3@��/���@        ��b:��*@��/���@        z�5��@���-��@        z�5��@��/���@        ��#�� @��/���@        ��#�� @��/����?                ��/����?        ��#�� @                        �cp>@        ��#��@                        �cp>@        ���>��@��/����?        ���>��@                        ��/����?        z�5��@                ��#���?                ;��,��@                        �cp>@        Ey�5A@��/���@        Dy�5A@��/����?        z�5��(@��/����?        ��#�� @                ��#��@��/����?        ��#��@                        ��/����?        �k(���5@                ��#���?                <��,��4@                        �cp>@                ��/����?                ��/����?        �k(��2@��/���.@0#0# @;��,��@��On�(@        ;��,��@��/���@        ��#��@��/����?                ��/����?        ��#��@                ��#���?�cp>@        ��#���?                        �cp>@                D�JԮD!@                �cp>@                �cp>@        ��b:��*@�cp>@0#0# @��#���?�cp>@        ��#���?                        �cp>@        z�5��(@        0#0# @<��,��$@                ��#�� @        0#0# @                0#0# @��#�� @                z�5��@�cp>'@        z�5��@��/���@                ��/���@        z�5��@                        ��/���@        Dy�5A@��/����?0#0#�?��#��@@��/����?        z�5��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ��#��@                ��b:��:@                ��#���?        0#0#�?                0#0#�?��#���?                �#���9@                z�5��@E�JԮD1@�C=�C=@                0#0#@z�5��@E�JԮD1@H�4H�4@��#���?                ��#�� @D�JԮD1@H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@��#�� @��/���.@                E�JԮD!@        ��#�� @���-��@                ���-��@        ��#�� @                ��b:��*@=l��F:B@0#0#�?��#�� @F�JԮDA@                0����/#@        ��#�� @��On�8@        ��#��@��On�8@        ��#�� @                ��#�� @��On�8@                ��On�(@        ��#�� @��On�(@        ��#���?                ��#���?��On�(@        ��#���?�cp>@                �cp>@        ��#���?                        0����/#@                ��/����?                ��/���@        ��#��@                ��#�� @                ��#�� @                ;��,��@��/����?0#0#�?��#��@                ��#���?��/����?0#0#�?��#���?        0#0#�?                0#0#�?��#���?                        ��/����?        �,����7@���-��:@)S2%S2G@�,����7@���-��:@�C=�C=<@�k(���5@h
��6@H�4H�4(@        �cp>'@0#0# @        0����/@0#0# @        �cp>@0#0# @        �cp>@0#0# @                0#0# @        �cp>@                        H�4H�4@        ��/����?                ���-��@        �k(���5@鰑%@0#0#@;��,��$@                [Lg1��&@鰑%@0#0#@z�5��@鰑%@0#0#@z�5��@鰑%@0#0# @                0#0# @z�5��@鰑%@        ��#�� @E�JԮD!@                E�JԮD!@        ��#�� @                ��#��@��/����?        ��#��@                        ��/����?                        0#0# @;��,��@                ��#�� @0����/@0#0#0@��#�� @0����/@H�4H�4@        0����/@H�4H�4@        0����/@                        H�4H�4@��#�� @                                ��8��8*@                vb'vb'2@                H�4H�4@                �A�A.@��#�� @��/���.@6��-�rW@��#�� @                        ��/���.@3��-�rW@        ��/����?                ���-��*@2��-�rW@                ��+��+D@        ���-��*@������J@        ��/����?%S2%S27@        ��/����?0#0# @        ��/����?H�4H�4@        ��/����?                        H�4H�4@                ��+��+@                �A�A.@        ��On�(@�A�A>@        �cp>'@�A�A.@        �cp>@�C=�C=,@        �cp>@0#0# @        ��/����?                ��/����?0#0# @        ��/����?                        0#0# @        �cp>@H�4H�4(@                0#0# @        �cp>@0#0#@        ��/����?                ��/����?0#0#@        ��/����?0#0#�?        ��/����?                        0#0#�?                H�4H�4@        �cp>@0#0#�?        �cp>@                        0#0#�?        ��/����?�A�A.@                �A�A.@        ��/����?        �t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��(.hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK݅�h��BX0         �                 ���?ʚB�S�?'      ���7{}@                        �jx?��S�W��?�       r^��vy@       ^                 ���@?wJ���?�       -$c)��l@                          �G�?;0Y�7�?g       ���xe@                         �!�?�l��f�?       �3f��:@������������������������       �               ��#��@                        �vQ?4>櫐�?       ��j���6@                         `<��?b%@�"�?       �6�E�1@	       
                  �6�?�����?       �O��@������������������������       �               ��/����?������������������������       �               ;��,��@                        8s�v? �F���?       :�.�-'@                       ���I?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �      �<       ��/���@                        \սP?      �<       0����/@������������������������       �               ��/����?������������������������       �               �cp>@       #                 �@�?��=r��?V       ='�[�a@                        �<��>�uE�~q�?       �ʷ��B@                        ��p?���/��?       V��7�@������������������������       �               ��/���@������������������������       �               ��#��@       "                 q��?Pdv���?       �2���=@                        0��?�]���?       �j0�W�<@                           �?��#�Ѵ�?       �)�B�4@������������������������       �        
       ��,���1@                        ��5?dn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @        !                 `��?�����?       ��X�)B @������������������������       �               ��/����?������������������������       �      ��       z�5��@������������������������       �               0#0#�?$       ?                 ��?��_;�*�?@       �si�A�Y@%       :                 �U���������?"       Lnj$O@&       9                 0fL�?����B�?       V=c$3 ?@'       ,                 �Ԏ?6�����?       �^��=@(       )                 �I?$ k�Lj�?       �q��l}@������������������������       �               ��/����?*       +                 ���s?`%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?-       8                    �?`n����?       � ��w<8@.       7                 �K��?��U�?        {|37@/       2                 0��?�_�A�?       ."�=LH5@0       1                 `��u?
4=�%�?       �(J��@������������������������       �               ��#�� @������������������������       �               �cp>@3       6                 ��?NF�X��?       .�=k�U0@4       5                 �:y?J9�)\e�?       _���b @������������������������       �               ;��,��@������������������������       �               �cp>@������������������������       �      ��       ��#�� @������������������������       �      м       ��/����?������������������������       �               ��#���?������������������������       �               0#0# @;       <                 ����?�	�� ��?       A�x��>@������������������������       �               ZLg1��6@=       >                 ���?��6L�n�?       �E#��h @������������������������       �               ��/����?������������������������       �      �<       ���>��@@       [                  ��?E���w��?       o�df_�D@A       H                 @�r�?C1����?       �/��l�A@B       E                 �_?�?�4�fP�?       V���-@C       D                  L��?�+�z���?	       KGh��
)@������������������������       �               0#0#�?������������������������       �      ��       �cp>'@F       G                 |�L?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?I       Z                 @��?k<S>	�?       S܃���4@J       U                  ���?;������?       �{f6�0@K       T                 �H��?�!�GU�?       m�����%@L       S                 �[�Z?LH����?       ��ϭ
*@M       R                 Эi�?|�G���?       ��%�|@N       O                 �!��?|��`p��?       �����@������������������������       �               0#0#�?P       Q                 ����?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               z�5��@������������������������       �      м       ��/���@V       Y                 �?��?��]ۀ��?       E���O@W       X                 �2�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               0#0#@������������������������       �               0#0#@\       ]                 �j%?      �<       z�5��@������������������������       �               ;��,��@������������������������       �               ��#���?_       x                 ��+a?<�)"(�?)       m�<99O@`       e                  @mj�?��,Yj�?#       9$���IK@a       b                 ��9�?�c�_��?       �/��=@������������������������       �               �cp>�9@c       d                    �?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@f       s                   p��?F�<�z�?       �7��S�8@g       r                 ���O?^�Jm�?       ��E�ǹ4@h       i                   �P�?trqw�H�?       i��Ч2@������������������������       �               ��#�� @j       o                 0��? +u�T�?       KDJ�ٕ0@k       l                 (��`?�}	;	�?	       vK�>4%@������������������������       �               0#0#�?m       n                 �5��>      �<       /����/#@������������������������       �               ��/����?������������������������       �               D�JԮD!@p       q                 ����?���/��?       @z$S��@������������������������       �               z�5��@������������������������       �               �cp>@������������������������       �      ܼ       ��#�� @t       u                 �C�P?f,���O�?       ���/>@������������������������       �               0#0# @v       w                  ��g�?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?y       z                  P(B�?|�G���?       ��%�|@������������������������       �               �cp>@{       ~                  `%+�?�@����?       ���a�@|       }                    �?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       H�4H�4@�       �                 ��0}?��ϵ��?k       Řﯞf@�       �                 �z?��2(&�?       �e4��\.@�       �                 �x�y?�D#���?       �B�j@������������������������       �               0#0#@������������������������       �               ��#�� @������������������������       �               vb'vb'"@�       �                 0��?�RZj�?c       hR|��3d@�       �                 �$�c?D��8�#�?(       ���1�3P@�       �                 P #�?����=��?       ���\?�H@�       �                  ��9?D�H���?       �S�m��G@�       �                 �=l�?Bǵ3���?       �q�ͨ�@������������������������       �               z�5��@�       �                 pH�?      �<       0����/@������������������������       �               ��/����?������������������������       �               ��/���@�       �                 @�?^���\�?       �E�S2�C@������������������������       �        	       ��b:��*@�       �                 �ګ?�S��W��?       $$�
�g:@������������������������       �               ��/����?�       �                 ����?�<�Aw��?       8&�+o|8@�       �                 XFe�?JH����?       ��ϭ
*@������������������������       �               z�5��@�       �                 ����?|�G���?       ��%�|@������������������������       �               ��/����?�       �                 �~N?|��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?�       �                 `U�?�x�<�?
       X&b��q1@�       �                 8vb�?      �<       z�5��(@������������������������       �               ��#���?������������������������       �               [Lg1��&@�       �                  A�?ޗZ�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@�       �                 �$ȧ?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?�       �                    �?      �<	       �A�A.@������������������������       �               vb'vb'"@������������������������       �               H�4H�4@�       �                 �6SZ?J� P��?;       �6��3X@�       �                 pHF�?x-�	X��?       n]�@��H@�       �                  �P�?�y�	��?       �Ͼ�w>@�       �                 ��0�?�4�fP�?
       X���-@������������������������       �               ���-��@�       �                 ѻ�?3y�d��?       �)h�2@�       �                 ���?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?�       �                 x��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/���@�       �                 h��?h/&$�S�?
       ���:�/@�       �                  ���?������?       +x�1�)@�       �                 �Ò=?\����?       Q	K��@������������������������       �      �<       z�5��@������������������������       �      ȼ       ��/����?������������������������       �               �cp>@������������������������       �               H�4H�4@������������������������       �      ��       /����/3@�       �                 ��O�?|�Ld�?       F����G@�       �                 ��I�?�'z�3�?       ���da�%@�       �                  0B�?���mf�?       寠�?b@������������������������       �      ��       ��/���@������������������������       �               0#0#�?������������������������       �               H�4H�4@�       �                 �1a�? ʊs`�?       �	S\!B@�       �                 p���?      �<       dJ�dJ�A@������������������������       �               0#0#�?������������������������       �               S2%S2%A@������������������������       �      �<       ��/����?�       �                 Б0�?�U�6�?,       rP)]P@�       �                  �Ԧ�?��弼�?)       �	x�p�N@�       �                 Фͽ?a{���?       �~8�31@������������������������       �               �cp>@�       �                 ����?vN��_�?       X��L,@�       �                 �N��?J5�,�r�?       7�r|k\@�       �                 TSK?����|e�?       �z �B�@������������������������       �               0#0# @�       �               ��~3�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               z�5��@�       �                  �u��?      �<       �C=�C=@������������������������       �               0#0#�?������������������������       �               H�4H�4@�       �                 0�Ь?��К���?       k�[��)F@�       �                 ��1�?Hy��]0�?       ���y"@������������������������       �               ��/����?������������������������       �               ��+��+@������������������������       �      ��       ��)��)C@�       �                  X3�?$�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?�t�bh�hhK ��h��R�(KK�KK��h �B�  ���khc@�B�)Dd@�؉��Ic@U^Cyc@�JԮDmc@f'vb'�X@��b:��Z@��On�X@%S2%S27@~�5��X@]�v%jWK@�C=�C=,@;��,��$@Nn��O0@        ��#��@                z�5��@Nn��O0@        z�5��@�cp>'@        ;��,��@��/����?                ��/����?        ;��,��@                ��#���?鰑%@        ��#���?�cp>@        ��#���?                        �cp>@                ��/���@                0����/@                ��/����?                �cp>@        �GpAV@1����/C@�C=�C=,@Ip�}>@���-��@0#0#�?��#��@��/���@                ��/���@        ��#��@                �#���9@�cp>@0#0#�?
�#���9@�cp>@        ������3@��/����?        ��,���1@                ��#�� @��/����?                ��/����?        ��#�� @                z�5��@��/����?                ��/����?        z�5��@                                0#0#�?    �M@�]�ڕ�?@��8��8*@�,����G@��On�(@0#0# @��,���1@�cp>'@0#0# @��,���1@�cp>'@        ��#���?��/���@                ��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#��0@��/���@        �P^Cy/@��/���@        �P^Cy/@�cp>@        ��#�� @�cp>@        ��#�� @                        �cp>@        ��b:��*@�cp>@        ;��,��@�cp>@        ;��,��@                        �cp>@        ��#�� @                        ��/����?        ��#���?                                0#0# @Kp�}>@��/����?        ZLg1��6@                ���>��@��/����?                ��/����?        ���>��@                [Lg1��&@1����/3@#0#0&@;��,��@1����/3@#0#0&@��#���?��On�(@0#0#�?        �cp>'@0#0#�?                0#0#�?        �cp>'@        ��#���?��/����?        ��#���?                        ��/����?        ��#��@���-��@��+��+$@��#��@���-��@H�4H�4@z�5��@�cp>@0#0# @z�5��@��/����?0#0# @        ��/����?0#0# @        ��/����?0#0# @                0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?        z�5��@                        ��/���@        ��#���?��/����?0#0#@��#���?��/����?                ��/����?        ��#���?                                0#0#@                0#0#@z�5��@                ;��,��@                ��#���?                ��#�� @�'�xr�F@vb'vb'"@��#�� @�)�B�D@��+��+@        ��|��<@0#0#�?        �cp>�9@                �cp>@0#0#�?                0#0#�?        �cp>@        ��#�� @��On�(@0#0#@���>��@��On�(@0#0#�?;��,��@��On�(@0#0#�?��#�� @                z�5��@��On�(@0#0#�?        /����/#@0#0#�?                0#0#�?        /����/#@                ��/����?                D�JԮD!@        z�5��@�cp>@        z�5��@                        �cp>@        ��#�� @                ��#���?        H�4H�4@                0#0# @��#���?        0#0#�?                0#0#�?��#���?                        ��/���@0#0#@        �cp>@                ��/����?0#0#@        ��/����?0#0#�?        ��/����?                        0#0#�?                H�4H�4@�GpAF@�a#6�K@��)��)S@��#�� @        ��8��8*@��#�� @        0#0#@                0#0#@��#�� @                                vb'vb'"@���#8E@�a#6�K@T��N��O@��,���A@��On�(@S2%S2%1@��,���A@��On�(@0#0# @��,���A@鰑%@0#0# @z�5��@0����/@        z�5��@                        0����/@                ��/����?                ��/���@        ���b:@@�cp>@0#0# @��b:��*@                �k(��2@�cp>@0#0# @        ��/����?        �k(��2@��/���@0#0# @z�5��@��/����?0#0# @z�5��@                        ��/����?0#0# @        ��/����?                ��/����?0#0# @                0#0# @        ��/����?        �P^Cy/@��/����?        z�5��(@                ��#���?                [Lg1��&@                z�5��@��/����?                ��/����?        z�5��@                        ��/����?                ��/����?                ��/����?                        �A�A.@                vb'vb'"@                H�4H�4@���>��@��]�ڕE@$S2%S2G@���>��@1����/C@0#0#@���>��@0����/3@0#0#@��#���?��On�(@0#0#�?        ���-��@        ��#���?�cp>@0#0#�?��#���?        0#0#�?��#���?                                0#0#�?        �cp>@                ��/����?                ��/���@        z�5��@���-��@H�4H�4@z�5��@���-��@        z�5��@��/����?        z�5��@                        ��/����?                �cp>@                        H�4H�4@        /����/3@                0����/@��-��-E@        ��/���@�C=�C=@        ��/���@0#0#�?        ��/���@                        0#0#�?                H�4H�4@        ��/����?dJ�dJ�A@                dJ�dJ�A@                0#0#�?                S2%S2%A@        ��/����?        z�5��@���-��@�;�;K@z�5��@0����/@������J@z�5��@��/���@��+��+$@        �cp>@        z�5��@��/����?��+��+$@z�5��@��/����?H�4H�4@        ��/����?H�4H�4@                0#0# @        ��/����?0#0#�?                0#0#�?        ��/����?        z�5��@                                �C=�C=@                0#0#�?                H�4H�4@        ��/����?�
��
�E@        ��/����?��+��+@        ��/����?                        ��+��+@                ��)��)C@        ��/����?0#0#�?        ��/����?                        0#0#�?�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJx�+hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK���h��B�5         �                  ����?����?�?,      ���T�}@       m                 ��ا?��=u'��?�       �>b2"wq@       *                 ���s?$"�i��?�       ����Bj@       #                 ��]"?�������?1       �W��'S@       "                 �p�?�17��?       ��r<�F@                        H��>���/��?       ��(�D@                        @��>~�����?       �4^$4�#@������������������������       �               ��#�� @	                        0?p�r{��?       e�6� @
                        ����?ʔfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               ��/���@                        "?�A&w(�?       �]��@@������������������������       �               ���>��@                        pTF�?p�Y�`��?       �����8@                         �\�?J�����?       g�C���3@                         ��n?d�r{��?       e�6� @������������������������       �               ���-��@������������������������       �               ��#���?                        @�E?���/��?       @z$S��'@                        ���U?�����?       ��X�)B @                        �-�?f%@�"�?       ��[�@������������������������       �               ��/����?                         �3��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ��       ;��,��@������������������������       �      ��       ��/���@       !                 Њ�(?�d�$���?       �T�f@                          h��?����?       ��X�)B@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?������������������������       �               ��#���?������������������������       �      �       ��/���@$       '                 �C>?k� ѽ?       �����>@%       &                 @��>`7uV��?        m}�'�:@������������������������       �               ��/����?������������������������       �      ��       �#���9@(       )                 p��A?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@+       \                 �6�?H�D�;�?T       �o:���`@,       U                 ��?}* 2N��??       �UΔKY@-       J                 �
o?g0�S��?2       {"�(iT@.       /                   ��?\ۀ]~��?        ̈�:K@������������������������       �               ��On�(@0       ?                 �U��><4��<�?       ��VS��D@1       2                 `Fe�?$_���1�?       d�&v�8@������������������������       �               ��#��@3       <                 �rQ�?Yf#�r�?       $(+m+�4@4       ;                  �P��?.�Cx@��?	       X�k�30@5       6                 ���Y?�=��	�?       .g�HH$@������������������������       �               ��/����?7       8                  @��?�wV����?       Bi�i�"@������������������������       �               ��#��@9       :                 -��?L� P?)�?       ����x�@������������������������       �               0#0#�?������������������������       �               ��#��@������������������������       �      Լ       �cp>@=       >                    �?      �<       0����/@������������������������       �               ��/���@������������������������       �               ��/����?@       A                 I#d?�(�����?
       ��0��0@������������������������       �               ��#�� @B       C                    �?l���A�?       0gX\-@������������������������       �               �cp>@D       I                 @F�fQ��?       �s�=�!@E       F                 � �?h%@�"�?       ��[�@������������������������       �               �cp>@G       H                 p茡?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      ��       �cp>@K       L                  p%+�?�D�+�?       Tx�-�;@������������������������       �               ��/����?M       P                 ��	�?.cÌ�v�?       `�u"��:@N       O                 �i�q?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?Q       T                 ����?8�u���?       ���i�7@R       S                 0kL�?�(1k��?       �ꁞ9�6@������������������������       �               �k(���5@������������������������       �      �<       ��/����?������������������������       �               0#0#�?V       W                 0*tC?�U1��-�?       8�KY��3@������������������������       �      ��	       �P^Cy/@X       [                 �^1�?�3`���?       .�r��@Y       Z                 k۬?���`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               ��#���?]       b                   ��?(s>.�?       �?�#@@^       _                 ��6�?�h��%�?
       �1�
�u0@������������������������       �      ��       ��|��,@`       a                 ����?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?c       l                 ���?F���u��?       ���KH�/@d       k                 P�$�?Ә�?ʊ�?
       ��l���)@e       f                ���${?l��w��?       ���@������������������������       �               ��/���@g       j                    �?�D#���?       �B�j@h       i                @u�2�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               0#0#�?������������������������       �               H�4H�4@������������������������       �      �<       �cp>@n       y                 0�2�?2�����?,       ����HWQ@o       p                 �#�?ܷB" �?       ���<�!:@������������������������       �               ��#��@q       x                  �~��?��H�&p�?       L^�3��5@r       w                 �/{�?hutee�?       P9��#@s       t                 0�!�?���mf�?       寠�?b@������������������������       �               �cp>@u       v                `�'�?v�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       ��+��+@������������������������       �               H�4H�4(@z       �                 j���?�������?       T����E@{       �                 �X\�?�F�g��?       �V���A@|       �                 �z>�?p̘�{7�?       �2}��]>@}       �                 �jE?����A�?       ��]���/@~       �                 ��>?As.�ʴ�?        E&A3*@       �                 ��|�?C��NV=�?       �t�ܲ@�       �                 @���?f%@�"�?       ��[�@������������������������       �               �cp>@�       �                 �R��?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               0#0# @������������������������       �      �<       ;��,��@������������������������       �      ��       �cp>@�       �                 |��?(�DNpk�?	       �k�Z$�,@�       �                 p���?,�b���?       �GXvƒ@������������������������       �               ;��,��@�       �                 ��V�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ���>��@������������������������       �      �       0����/@������������������������       �               0#0# @�       �                 oք?���~��?{       �Q�D�%h@�       �                 7b?�NP��R�?        �]���J@�       �                 eni?��j ��?       ��"�G@�       �                 �$'.?�0�0���?       ���ȐsC@�       �                 �y���B�A ��?       Bb�1�O8@�       �                 ����?�`@s'��?       Ei_y,*@������������������������       �               ��#���?������������������������       �               �cp>@�       �                 �?P�:V��?       �GP�1@�       �                  0���?����?       ��X�)B@�       �                 ��f?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �               ��b:��*@�       �                  `<��?��Ik���?	       ��c��.-@�       �                 �闾?lSmd�d�?       :��P{�@�       �                    �?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?�       �                    �?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ��       ���-��@�       �                 `Fe�?��t1u�?       "�te!� @������������������������       �               0#0#�?������������������������       �      ��       ���>��@������������������������       �               H�4H�4@�       �                 p'v�?~}����?[       W: �a@�       �                 �-4�?���[�k�?       �!�c�B@�       �                  f&�?,��V�"�?       ��y���/@�       �                 ��u�?�N�+�?	       ����*@�       �                 ����?�AP�9��?       i��6��@������������������������       �               ��+��+@������������������������       �      �<       ��/����?������������������������       �      ��       H�4H�4@�       �                 �(��?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                  P�?�˒�0�?       �A��Z!5@������������������������       �               �C=�C=,@�       �                  ���?d�ih�<�?       ��
@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                 @�/�?�N�y1��?C       ��/���Y@�       �                  ^M�?P1�+��?0       ^ܦGV.S@�       �                 �7�?��$eq��?       <���.C@�       �                 ��a�?�Yi�e?�?       ��3���8@�       �                 ��f?��M��,�?	       x��r�0@�       �                 �؉�?���#��?       Y�f���'@�       �                 P��?��[����?       Hl�_A@������������������������       �               0����/@������������������������       �               0#0# @�       �                 @	+�?�Z�	7�?       j~���@������������������������       �               ��/����?�       �                  �P�?�����?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?������������������������       �               0����/@�       �                 �0�?l�z���?       p���f @�       �                    �?f,���O�?       ���/>@�       �                 @o4�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               0#0# @������������������������       �               ��#��@�       �                 ��6�?�;�a
=�?	       ��l��+@������������������������       �      ��       鰑%@�       �                 ����?z��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?�       �                 �A�?4$��(�?       {����-C@�       �                 `Fe�?i=��?       *����%A@�       �                 pwG�?     ��?       "F�b@������������������������       �               H�4H�4@������������������������       �               ��#�� @�       �                 �fQ?P����D�?       ���2=@������������������������       �      ��       0#0#0@�       �                  �nY?�n���k�?       3��&�*@������������������������       �               ��/����?������������������������       �               H�4H�4(@�       �                 ���?
����?       ��X�)B@������������������������       �               ��#�� @�       �                 �у�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                    �?��}�d�?       �1$�~&:@�       �                 @8��?1����?       �`O��"@�       �                 uK�b?�`�ox��?       
c��0 @������������������������       �               ��#���?�       �                 TQQ�?      �<       �C=�C=@������������������������       �               0#0#�?������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?�       �                 P��?�6��b�?       %�|�1@�       �                 �؈�?�v�;B��?       ՟���	 @�       �                 P�$�?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               ��+��+@������������������������       �               vb'vb'"@�t�bh�hhK ��h��R�(KK�KK��h �B�  �#����e@鰑Nc@k�i��a@�5�װ`@��F:l$Z@�ڬ�ڬD@�>��n[@h
��V@H�4H�4(@�}�\I@�cp>�9@        �k(���5@�e�_��7@        �k(���5@'jW�v%4@        z�5��@���-��@        ��#�� @                ��#���?���-��@        ��#���?�cp>@                �cp>@        ��#���?                        ��/���@        �k(��2@���-��*@        ���>��@                \Lg1��&@���-��*@        ���>��@��On�(@        ��#���?���-��@                ���-��@        ��#���?                z�5��@�cp>@        z�5��@��/����?        ��#���?��/����?                ��/����?        ��#���?��/����?        ��#���?                        ��/����?        ;��,��@                        ��/���@        ��#��@��/����?        z�5��@��/����?        z�5��@                        ��/����?        ��#���?                        ��/���@        ���>��<@��/����?        �#���9@��/����?                ��/����?        �#���9@                z�5��@��/����?                ��/����?        z�5��@                    �M@1����-O@H�4H�4(@,�����K@�)�B�D@0#0#@������C@&jW�v%D@0#0# @��#��0@;l��F:B@0#0#�?        ��On�(@        ��#��0@�e�_��7@0#0#�?z�5��(@�cp>'@0#0#�?��#��@                ��#�� @�cp>'@0#0#�?��#�� @���-��@0#0#�?��#�� @��/����?0#0#�?        ��/����?        ��#�� @        0#0#�?��#��@                ��#��@        0#0#�?                0#0#�?��#��@                        �cp>@                0����/@                ��/���@                ��/����?        ��#��@��On�(@        ��#�� @                ��#�� @��On�(@                �cp>@        ��#�� @���-��@        ��#�� @��/���@                �cp>@        ��#�� @��/����?        ��#�� @                        ��/����?                �cp>@        \Lg1��6@��/���@0#0#�?        ��/����?        \Lg1��6@�cp>@0#0#�?��#���?��/����?        ��#���?                        ��/����?        �k(���5@��/����?0#0#�?�k(���5@��/����?        �k(���5@                        ��/����?                        0#0#�?��#��0@��/����?0#0# @�P^Cy/@                ��#���?��/����?0#0# @        ��/����?0#0# @                0#0# @        ��/����?        ��#���?                z�5��@鰑5@0#0# @��#�� @��|��,@                ��|��,@        ��#�� @                ��#���?                ��#���?                ��#���?���-��@0#0# @��#���?��/���@0#0# @��#���?��/���@0#0# @        ��/���@        ��#���?        0#0# @��#���?        0#0#�?��#���?                                0#0#�?                0#0#�?                H�4H�4@        �cp>@        �,����7@Nn��O0@�s?�s?=@��#��@��/���@vb'vb'2@��#��@                        ��/���@vb'vb'2@        ��/���@H�4H�4@        ��/���@0#0#�?        �cp>@                ��/����?0#0#�?        ��/����?                        0#0#�?                ��+��+@                H�4H�4(@������3@��On�(@#0#0&@������3@��On�(@H�4H�4@������3@��/���@H�4H�4@���>��@���-��@0#0# @���>��@��/���@0#0# @��#�� @��/���@0#0# @��#�� @��/���@                �cp>@        ��#�� @��/����?                ��/����?        ��#�� @                                0#0# @;��,��@                        �cp>@        z�5��(@��/����?0#0#�?;��,��@��/����?0#0#�?;��,��@                        ��/����?0#0#�?        ��/����?                        0#0#�?���>��@                        0����/@                        0#0# @���#8E@��On�H@r�6k�6Y@��b:��:@:l��F:2@0#0# @��b:��:@;l��F:2@0#0# @������3@:l��F:2@0#0#�?��,���1@���-��@        ��#���?�cp>@        ��#���?                        �cp>@        ��#��0@��/����?        z�5��@��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#�� @                ��b:��*@                ��#�� @�cp>'@0#0#�?��#�� @0����/@0#0#�?        �cp>@0#0#�?        �cp>@                        0#0#�?��#�� @��/����?                ��/����?        ��#�� @                        ���-��@        ���>��@        0#0#�?                0#0#�?���>��@                                H�4H�4@�P^Cy/@�]�ڕ�?@+S2%S2W@��#���?0����/@=�C=�C?@��#���?��/���@#0#0&@        ��/����?#0#0&@        ��/����?��+��+@                ��+��+@        ��/����?                        H�4H�4@��#���?��/����?        ��#���?                        ��/����?                ��/����?��+��+4@                �C=�C=,@        ��/����?H�4H�4@        ��/����?                        H�4H�4@���>��,@���-��:@0��+��N@��b:��*@��On�8@��)��)C@��#�� @�cp>7@�C=�C=@��#�� @�cp>'@��+��+@z�5��@�cp>'@0#0# @z�5��@���-��@0#0# @        0����/@0#0# @        0����/@                        0#0# @z�5��@��/����?                ��/����?        z�5��@��/����?        z�5��@                        ��/����?                0����/@        ;��,��@        H�4H�4@��#���?        H�4H�4@��#���?        0#0#�?��#���?                                0#0#�?                0#0# @��#��@                        �cp>'@0#0# @        鰑%@                ��/����?0#0# @                0#0# @        ��/����?        ;��,��@��/����?=�C=�C?@��#�� @��/����?=�C=�C?@��#�� @        H�4H�4@                H�4H�4@��#�� @                        ��/����?�C=�C=<@                0#0#0@        ��/����?H�4H�4(@        ��/����?                        H�4H�4(@z�5��@��/����?        ��#�� @                ��#���?��/����?        ��#���?                        ��/����?        ��#���?��/����?%S2%S27@��#���?��/����?�C=�C=@��#���?        �C=�C=@��#���?                                �C=�C=@                0#0#�?                H�4H�4@        ��/����?                ��/����?0#0#0@        ��/����?�C=�C=@        ��/����?0#0# @        ��/����?                        0#0# @                ��+��+@                vb'vb'"@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJH�SshFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKх�h��B�-         �                 p��g?0�U��#�?6      �(��}@       �                 `m�?p����?�       b���-wv@       �                 (/��?0�U�B6�?�       ����Hr@       S                    �?�]�R�?�       	IY��(r@                        P�hf?�1R��?r       pt'�/g@                        � C;?V*�"�?.       jܤ?[�S@                        �+"�?  	$�?)       ���*Q@       	                  �Ԧ�?\��e�)�?'       UVl��P@������������������������       �               �cp>@
                        �U���������?%       8nҟ��O@                         Q�J?`Տ�m|�?       ��h
�7@                        T�@?^n����?	       � ��w<(@                         �~��?ʔfm���?       ��Z�N@������������������������       �               ��/����?                          �P�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?                        �c-?|�6L�n�?       �E#��h @������������������������       �      �<       ���>��@������������������������       �      ȼ       ��/����?                        ���f?      �<       [Lg1��&@������������������������       �               ��#�� @������������������������       �               �k(��"@������������������������       �      ��       ��k(/D@������������������������       �      	�       ��/����?                        0��?������?       �4^$4�#@                       @* r?      �<       ���-��@������������������������       �               ��/���@������������������������       �               �cp>@������������������������       �               z�5��@       $                 ��{�?�x�'��?D       �DӿZ@        !                  ��d�?�@G���?       X��Q7@������������������������       �               ��On�(@"       #                 h3�?��Ñp��?       <7��0�%@������������������������       �               0����/@������������������������       �               H�4H�4@%       B                 �T�x?�Q�m��?6       2 �%_�T@&       9                 `�г?�\U�?       �{����G@'       6                 ��?��*F��?       j�;=�nA@(       +                 �E�?�����?       \��j>@)       *                 �;�?l@ȱ��?	       nm���S'@������������������������       �               ��#�� @������������������������       �      ��       /����/#@,       3                 px��?�����?	       L��o�g2@-       .                 �j%?^P�D�?       �A��P?$@������������������������       �               z�5��@/       2                 h�R?Ȕfm���?       ��Z�N@0       1                 ��[r?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��#���?4       5                 8X9�?      �<       ��#�� @������������������������       �               ��#�� @������������������������       �               z�5��@7       8                 \��?      �<       0����/@������������������������       �               ��/����?������������������������       �               ��/���@:       A                 P	��?u�Z\�?	       eA�F/*@;       <                 йu�?�K��t�?       N����"@������������������������       �               ��/����?=       >                  �jw?�.�KQu�?       �K̎@������������������������       �               ��#�� @?       @                 X�˙?�o���?       o�9�F@������������������������       �               0#0#@������������������������       �               ��#���?������������������������       �               0#0#@C       P                 `A��?�8u#��?       ��_O;�A@D       I                 ��g�?�w��?       ���4?_@@E       F                 ��?���P��?       �*Y�ȹ9@������������������������       �               ������3@G       H                 ��W�?hn����?       � ��w<@������������������������       �      ȼ       ��/����?������������������������       �               ��#��@J       O                 @�ĥ?�)z� ��?       ~�\�@K       N                 ��:�?Ĕfm���?       ��Z�N@L       M                 p��A?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               z�5��@Q       R                 8�]�?���`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @T       �                 `&�?�vU�T�?L       
D|�CZ@U       Z                 ��R?�T��V��?:       =cn��`T@V       Y                 ���k?`�s�	�?       e���*@W       X                 0Ŕ>?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               <��,��$@[       p                 ��?p������?2       �a�j|Q@\       ]                 ����?�5T501�?       �o8\�8@������������������������       �               ��#�� @^       i                 P�^�?2$ĝ��?       �P�3ew6@_       `                 8qL1?64|���?       	�T|qt2@������������������������       �               E�JԮD!@a       h                   ���?������?	       �4^$4�#@b       c                 �΢뾤��/��?       @z$S��@������������������������       �               ��/����?d       e                 @F�����?       ��X�)B@������������������������       �               ��#���?f       g                 8*��?bn����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      ��       ��/���@j       m                 �\�?�3`���?       .�r��@k       l                  E(�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?n       o                   �0�?      �<       0#0# @������������������������       �               0#0#�?������������������������       �               0#0#�?q       �                 @�?� �����?       �:�J�E@r       {                  �Є?RsaѠ�?       <�k(=@s       z                 �?�?���+���?       ���h�0@t       w                  P���? 3�Ҽ��?       ����@,@u       v                 P��x?*k�"O��?       �?<��*&@������������������������       �      ��       ���>��@������������������������       �      ȼ       ��/���@x       y                 ����?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �      �<       �cp>@|       }                 �u�?�����?	       �O��(@������������������������       �               ��/����?~                        �f�?����X��?       &��֞&@������������������������       �      ��       <��,��$@������������������������       �      ȼ       ��/����?�       �                 �S�?\Lj����?       ���T�,@������������������������       �               z�5��(@������������������������       �               0#0# @�       �                 ��f�?R��US��?       9�7���7@�       �                  h��?����|e�?       �z �B�@�       �                 0�"]?lutee�?       Q9��@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               H�4H�4@�       �                 p|߰?�	>�S�?       ���FV%/@�       �                 ��n�?�)��R=�?
       �
3�e1)@������������������������       �               ��#���?�       �                  0Y��?�>s{Ab�?	       aI��n'@������������������������       �               鰑%@������������������������       �               0#0#�?�       �                ��!�?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �     ��       0#0# @�       �                 j:?���̊�?)       kmh�۸P@�       �                 �vQ?����8V�?       ;�tB̢H@�       �                 �R�־��&���?       �p4���@@�       �                  v�?�P1���?        � ?@�       �                   �x�?��
+���?       \Zz�+�#@������������������������       �               0����/@�       �                 ���?L� P?)�?       ����x�@������������������������       �               ��#��@������������������������       �               0#0#�?������������������������       �               ��-��-5@������������������������       �      �<       ��#�� @�       �                 �u�?l[
�ݢ�?
       F_�Ș0@�       �                 ��ٻ?��6L�n�?       �E#��h @������������������������       �               ��#��@�       �                 ��b�?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@�       �                 �m�?x�G���?       ��%�|@������������������������       �               ��/����?�       �                 ��C�?|��`p��?       �����@������������������������       �               0#0#@������������������������       �      �<       ��/����?�       �                   p��?�`���6�?       .u��֝1@�       �                 0p^�?��Ik���?       ��c��.-@�       �                 �� �?��2uj�?
       j溕+@�       �                    �?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �      ȼ       �cp>'@������������������������       �      �<       ��#���?������������������������       �               H�4H�4@�       �                 �=�t?��oH��?M       `�QI��\@������������������������       �               ��#���?�       �                 p�?H�O�T��?L       :A�hya\@�       �                 �}�?��#���?       �͆�1�2@������������������������       �               ��/����?�       �                 h~��?Jy��]0�?       �N-ۙ2@�       �                 `Qt�?r����?
       Qz�i0@�       �                 �N�X?      �<       ��8��8*@������������������������       �               0#0# @������������������������       �               #0#0&@�       �                 �+�[?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                ���;�?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?�       �                 �K�n?�S&�Ƨ�??       č ���W@�       �                 8�h�?�Qk��?       ��Th!�@�       �                    �?h�4���?       �tCP��@������������������������       �               0#0#�?�       �                 Ќ�j?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �               0#0# @�       �                  �?���##�?:       g>��J�U@�       �                 �Q�?      �<.       zb'vb'R@������������������������       �               0#0# @������������������������       �        -       fJ�dJ�Q@�       �                 �s�?h�E�B��?       dߞKC.@������������������������       �               ��/����?������������������������       �               ��8��8*@�t�b�!     h�hhK ��h��R�(KK�KK��h �B�  �GpAf@��`@�fm�f�d@     f@s�����]@=�C=�CO@��k(/d@3�@S�X@0#0#@@��k(/d@0�@S�X@�A�A>@.�����[@��|��L@0#0#0@$�}��O@��/���.@        Kp�}N@D�JԮD!@        Lp�}N@���-��@                �cp>@        Mp�}N@��/���@        ������3@��/���@        ��#�� @��/���@        ��#���?�cp>@                ��/����?        ��#���?��/����?        ��#���?                        ��/����?        ���>��@��/����?        ���>��@                        ��/����?        [Lg1��&@                ��#�� @                �k(��"@                ��k(/D@                        ��/����?        z�5��@���-��@                ���-��@                ��/���@                �cp>@        z�5��@                4��tSH@鰑E@0#0#0@        E�JԮD1@H�4H�4@        ��On�(@                0����/@H�4H�4@        0����/@                        H�4H�4@5��tSH@��On�8@��+��+$@<��,��4@0����/3@0#0# @��,���1@E�JԮD1@        ��,���1@��On�(@        ��#�� @0����/#@        ��#�� @                        /����/#@        �P^Cy/@�cp>@        ���>��@�cp>@        z�5��@                ��#���?�cp>@                �cp>@                ��/����?                ��/����?        ��#���?                ��#�� @                ��#�� @                z�5��@                        0����/@                ��/����?                ��/���@        z�5��@��/����?0#0# @z�5��@��/����?0#0#@        ��/����?        z�5��@        0#0#@��#�� @                ��#���?        0#0#@                0#0#@��#���?                                0#0#@*�����;@�cp>@0#0# @,�����;@0����/@        �,����7@��/����?        ������3@                ��#��@��/����?                ��/����?        ��#��@                ��#��@�cp>@        ��#���?�cp>@                �cp>@                ��/����?                ��/����?        ��#���?                z�5��@                        ��/����?0#0# @        ��/����?                        0#0# @~�5��H@�)�B�D@�C=�C=,@5��tSH@�a#6�;@��+��+@z�5��(@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        <��,��$@                �YLg1B@���-��:@��+��+@z�5��@On��O0@0#0# @��#�� @                ��#��@On��O0@0#0# @z�5��@��/���.@                E�JԮD!@        z�5��@���-��@        z�5��@�cp>@                ��/����?        z�5��@��/����?        ��#���?                ��#�� @��/����?        ��#�� @                        ��/����?                ��/���@        ��#���?��/����?0#0# @��#���?��/����?                ��/����?        ��#���?                                0#0# @                0#0#�?                0#0#�?Kp�}>@鰑%@H�4H�4@��,���1@鰑%@0#0#�?���>��@E�JԮD!@0#0#�?���>��@�cp>@0#0#�?���>��@��/���@        ���>��@                        ��/���@                ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@        <��,��$@��/����?                ��/����?        <��,��$@��/����?        <��,��$@                        ��/����?        z�5��(@        0#0# @z�5��(@                                0#0# @��#���?���-��*@vb'vb'"@        ��/����?H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@                H�4H�4@��#���?�cp>'@H�4H�4@��#���?鰑%@0#0#�?��#���?                        鰑%@0#0#�?        鰑%@                        0#0#�?        ��/����?0#0# @        ��/����?                        0#0# @                0#0# @�P^Cy/@鰑5@�A�A>@��b:��*@0����/#@��8��8:@z�5��@0����/@#0#06@��#��@0����/@#0#06@��#��@0����/@0#0#�?        0����/@        ��#��@        0#0#�?��#��@                                0#0#�?                ��-��-5@��#�� @                ���>��@0����/@0#0#@���>��@��/����?        ��#��@                z�5��@��/����?                ��/����?        z�5��@                        ��/���@0#0#@        ��/����?                ��/����?0#0#@                0#0#@        ��/����?        ��#�� @�cp>'@0#0#@��#�� @�cp>'@0#0#�?��#���?�cp>'@0#0#�?��#���?        0#0#�?                0#0#�?��#���?                        �cp>'@        ��#���?                                H�4H�4@��#���?D�JԮD!@��8��8Z@��#���?                        D�JԮD!@��8��8Z@        ��/���@�A�A.@        ��/����?                �cp>@�A�A.@        ��/����?�A�A.@                ��8��8*@                0#0# @                #0#0&@        ��/����?0#0# @        ��/����?                        0#0# @        ��/����?                ��/����?                ��/����?                0����/@��
�pV@        �cp>@0#0#@        �cp>@0#0# @                0#0#�?        �cp>@0#0#�?                0#0#�?        �cp>@                        0#0# @        ��/����?�~��~nU@                zb'vb'R@                0#0# @                fJ�dJ�Q@        ��/����?��8��8*@        ��/����?                        ��8��8*@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�8�hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK���h��B�5         t                  �~��?�+�O�?.      A��w}@       _                 �ŗ�?�5u��i�?}       �4iИ�h@       L                 �㨤?��l�*�?h       ��[V�d@                        �w�m?$�2�K�?Q       �/^�`@                        ����?�4����?       �Ӯ���C@                         ���?��Ik���?       ��c��.=@                        @��)?������?       �N0gX1@       	                   ��?r@ȱ��?       om���S@������������������������       �               ��/���@
                        d1O�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               �cp>'@                         �3��?���#��?       X�f���'@                        ���?�|2N��?       �3K}@������������������������       �               z�5��@������������������������       �               0#0# @������������������������       �      ��       ���-��@                        p��e?���/��?       6��o��#@������������������������       �               �cp>@                        ��??�_�A�?       肵�e`@                         @?��?���/��?       V��7�@������������������������       �               ��/����?                         �a�?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               z�5��@       7                 �x�.?&��`�?;       ҟ@��.X@       2                 ���?���d�?       �)�r�L@       /                 P���?�K���x�?       �
3�e1I@       &                 ��ͅ?��;���?       ���6:&G@        !                 hl��?.�r?�?       �M�)#�;@������������������������       �      ȼ       �k(��2@"       #                 ��s?h�j���?       ���z"@������������������������       �               ��/����?$       %                 �/��?      �<       ��#�� @������������������������       �               ��#�� @������������������������       �               z�5��@'       (                 0=T�?޺W�w��?       �'DQm2@������������������������       �               0#0# @)       *                 8LSR?|�6L�n�?
       �E#��h0@������������������������       �               ��/����?+       .                 08��?(k� ѽ?	       �����.@,       -                 0I��?����?       ��X�)B@������������������������       �      ��       z�5��@������������������������       �      �<       ��/����?������������������������       �               \Lg1��&@0       1                  �9��?�J���?       ��*]Y@������������������������       �               ��#�� @������������������������       �               0#0# @3       6                     �?�_�A�?       肵�e`@4       5                 ���?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               z�5��@8       G                 �͋?������?       W/O�C@9       @                  `S��?. k�Lj�?       e*�}#<=@:       ;                  G8W?���/��?       V��7�@������������������������       �               �cp>@<       ?                  `s�?�d�$���?       �T�f@=       >                 D�{e?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               z�5��@A       F                 ��?�^�#΀�?       O�{��A5@B       E                 �Q�?��٤ݸ?       ��<5�84@C       D                 @F�Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �      ��       On��O0@������������������������       �      �<       ��#���?H       K                   \��?i,�V�?       8����$@I       J                 �6�?���/��?       @z$S��@������������������������       �               z�5��@������������������������       �               �cp>@������������������������       �               0#0#@M       N                  `s�?�%��̫�?       !'`�'=@������������������������       �               ��#���?O       ^                 0�/�?v1���?       �8���<@P       ]                 �*��?$����?        X�[�;@Q       Z                 �
�k?䱐3+>�?       �'�8�:@R       W                 �:��?$NU�w�?       ���6:&7@S       V                 ��դ?�G�<�J�?       T �24@T       U                  �9��?�;�a
=�?       ��l��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �        
       ���-��*@X       Y                 tM�D?j%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?[       \                    �?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �      �<       ��#���?`       s                 @Q�?��:m��?       +eª�?@a       b                 �$I�?ΗP����?       |t��"�:@������������������������       �               ��+��+@c       d                  "��?"��x1�?       ̓�L2�5@������������������������       �               0#0# @e       p                 0I��?������?       �#�ҏ3@f       i                 �X�?:ĩAf�?       ��d>v�0@g       h                �e:s�?�5JH���?       �MOI#@������������������������       �               E�JԮD!@������������������������       �               0#0#�?j       o                 �e_�?��|��?       ���ĺw@k       l                 @�t�?`n����?       � ��w<@������������������������       �               ��#���?m       n                 ��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       ��/���@q       r                 @}��?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               ��+��+@u       �                 �]�?��.d�:�?�       �4�h�+q@v       �                 ��\�?`��"/��?[       ;U6�b@w       �                 0׋w?��q�R�?L       ����rG]@x       �                 ���?��$7��?8       �OsΎsT@y       �                 @?J�}�~�?       �2O�6�C@z       �                 �&pX?�d�$���?       ;�)�T�A@{       �                 ����?�N,u��?       ��u�=@|       �                   ���?h�j���?       ^��\�;@}       ~                 ��V?��Z�	7�?       j~���@������������������������       �               ��#�� @       �                 ����?f%@�"�?       ��[�@������������������������       �               ��/����?�       �                 8/h?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 �y����(1k��?       �ꁞ9�6@�       �                 �k�J?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@������������������������       �      м       �k(��2@�       �                    �?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                  �?���/��?       Az$S��@������������������������       �               �cp>@�       �                 �3�_?      �<       z�5��@������������������������       �               ��#�� @������������������������       �               ��#���?�       �                  �!�?�fm���?       ��Z�N@�       �                 h��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 �\3�?����rk�?       |l��E@�       �                 P�Dv?v	����?        ��>�A@�       �                 @Ws�?�0�����?       ��Ʃ6@������������������������       �               H�4H�4@�       �                   �x�?�(�����?
       ��0��0@�       �                 �m�?�d�$���?       �T�f@������������������������       �               ��/����?�       �                 H��>      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@������������������������       �      Լ       �cp>'@������������������������       �               ��On�(@�       �                 l'��?      �<       �C=�C=@������������������������       �               0#0#�?������������������������       �               H�4H�4@�       �                 p��?�� M�?       �Q�4ȧA@�       �                  `s�?+�d���?       ��{h&@�       �                 0�2�?�����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?�       �                 (�i<?�o���?       o�9�F@������������������������       �               ��#���?������������������������       �               0#0#@�       �                 ��a?v=���?       � ��R8@�       �                 ��W9?|�G���?       ��%�|@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �        	       ��+��+4@�       �                 PWe|?�!:de�?       &�&ޔ�;@�       �                 �Ua'?���/��?       6��o��#@�       �                 ���?��|��?       ���ĺw@�       �                 h���?^n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               ��/���@�       �                  �6��?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �        
       ��,���1@�       �                 ����?NII{���?V       ����A`@�       �                  ����?~T�#q�?)       �&qP@�       �                  jZ?�=
���?(       �G�N@�       �                 �W�?���o:��?       ��l���=@������������������������       �               �cp>@�       �                 ��Ĳ?�I�?       �%`/��:@�       �                 @��?pO6�?       �d�*ę8@�       �                 `��B?���o�:�?
       ����+@�       �                 p�?�]
���?       ��Ј�'@�       �                 �{��?޾�R���?       :�S) $@�       �                  ���?:�N9���?       ��{j�@������������������������       �               ��/����?�       �                 pEʦ?b,���O�?       ���/>@������������������������       �               ��#���?������������������������       �               H�4H�4@������������������������       �               ��+��+@������������������������       �      ȼ       ��/����?������������������������       �      м       ��/����?�       �                 @��?������?       +�ǟf%@�       �                 `ec�?����|e�?       �z �B�@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?������������������������       �               ���-��@������������������������       �      ܼ       ��#�� @�       �                 �Z�?�v�;B��?       ՟���	@@������������������������       �      ��       #0#06@�       �                 `�?�?putee�?       Q9��#@�       �                 ܆�?`�ih�<�?       ��
@�       �                  ���?|��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               0#0#@������������������������       �               �cp>@������������������������       �      �<       ��#��@�       �                 p���?HU�6�?-       tP)]P@�       �                  �rm?d�����?(       ���dߞL@�       �                 �dY�?�E���?       �|����4@�       �                 ,�u�?�� ��?       rp� k@�       �                  ���?���mf�?       寠�?b@�       �                 �<M�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �      ��       �cp>@������������������������       �               0#0#�?�       �                 �D����(v��?       �A�s(.@�       �                 ���?�v�;B��?       ՟���	 @������������������������       �               ��/����?������������������������       �               �C=�C=@������������������������       �               �C=�C=@�       �                ��5p�?      �<       vb'vb'B@������������������������       �               H�4H�4@������������������������       �               B�A�@@�       �                 x��?QH����?       ��ϭ
*@�       �                   ���?��Z�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@������������������������       �               0#0# @�t�bh�hhK ��h��R�(KK�KK��h �B�  ��Gp_b@��-��bd@��+��+d@��Gp_R@=�cp�W@�C=�C=<@��,���Q@��-��bT@��8��8*@"�}��P@G�)�BM@��+��+$@�k(��"@�a#6�;@0#0# @��#��@�cp>7@0#0# @��#���?On��O0@        ��#���?0����/@                ��/���@        ��#���?��/����?                ��/����?        ��#���?                        �cp>'@        z�5��@���-��@0#0# @z�5��@        0#0# @z�5��@                                0#0# @        ���-��@        ;��,��@0����/@                �cp>@        ;��,��@��/����?        ��#�� @��/����?                ��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        z�5��@                ���>��L@��/���>@0#0# @5��tSH@0����/@0#0#@�k(���E@�cp>@0#0#@=��,��D@�cp>@0#0# @��b:��:@��/����?        �k(��2@                ��#�� @��/����?                ��/����?        ��#�� @                ��#�� @                z�5��@                ���>��,@��/����?0#0# @                0#0# @���>��,@��/����?                ��/����?        ���>��,@��/����?        z�5��@��/����?        z�5��@                        ��/����?        \Lg1��&@                ��#�� @        0#0# @��#�� @                                0#0# @;��,��@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                z�5��@                �k(��"@�cp>�9@0#0#@z�5��@�cp>7@        ��#��@��/���@                �cp>@        ��#��@��/����?        ��#���?��/����?                ��/����?        ��#���?                z�5��@                ��#�� @/����/3@        ��#���?0����/3@        ��#���?�cp>@                �cp>@        ��#���?                        On��O0@        ��#���?                z�5��@�cp>@0#0#@z�5��@�cp>@        z�5��@                        �cp>@                        0#0#@z�5��@�cp>7@H�4H�4@��#���?                ��#�� @�cp>7@H�4H�4@��#���?�cp>7@H�4H�4@��#���?�cp>7@0#0# @��#���?鰑5@0#0#�?        1����/3@0#0#�?        �cp>@0#0#�?        �cp>@                        0#0#�?        ���-��*@        ��#���?��/����?        ��#���?                        ��/����?                ��/����?0#0#�?                0#0#�?        ��/����?                        0#0#�?��#���?                z�5��@���-��*@�A�A.@z�5��@���-��*@��+��+$@                ��+��+@z�5��@���-��*@��+��+@                0#0# @z�5��@���-��*@H�4H�4@��#�� @���-��*@0#0#�?        E�JԮD!@0#0#�?        E�JԮD!@                        0#0#�?��#�� @0����/@        ��#�� @��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                        ��/���@        ��#���?        0#0# @��#���?                                0#0# @                ��+��+@��Gp_R@��t�HQ@F�A�`@%�}��O@鰑E@������C@��k(/D@�+Q��B@������C@Fy�5A@F�JԮDA@��8��8*@Lp�}>@/����/#@        ���>��<@���-��@        �#���9@��/���@        |�5��8@�cp>@        z�5��@��/����?        ��#�� @                ��#���?��/����?                ��/����?        ��#���?��/����?                ��/����?        ��#���?                �k(���5@��/����?        z�5��@��/����?                ��/����?        z�5��@                �k(��2@                ��#���?��/����?        ��#���?                        ��/����?        z�5��@�cp>@                �cp>@        z�5��@                ��#�� @                ��#���?                ��#���?�cp>@                �cp>@                ��/����?                ��/����?        ��#���?                ��#��@��On�8@��8��8*@��#��@��On�8@H�4H�4@��#��@��On�(@H�4H�4@                H�4H�4@��#��@��On�(@        ��#��@��/����?                ��/����?        ��#��@                ��#���?                z�5��@                        �cp>'@                ��On�(@                        �C=�C=@                0#0#�?                H�4H�4@z�5��@�cp>@��8��8:@z�5��@��/����?0#0#@;��,��@��/����?        ;��,��@                        ��/����?        ��#���?        0#0#@��#���?                                0#0#@        ��/����?#0#06@        ��/����?0#0# @                0#0# @        ��/����?                        ��+��+4@ZLg1��6@0����/@        ;��,��@0����/@        ��#�� @0����/@        ��#�� @��/����?                ��/����?        ��#�� @                        ��/���@        z�5��@                ��#���?                ��#�� @                ��,���1@                ;��,��$@�cp>�9@6��-�rW@���>��@0����/3@������C@z�5��@1����/3@������C@z�5��@��/���.@#0#0&@        �cp>@        z�5��@��On�(@#0#0&@��#���?��On�(@#0#0&@��#���?0����/@0#0# @��#���?�cp>@0#0# @��#���?��/����?0#0# @��#���?��/����?H�4H�4@        ��/����?        ��#���?        H�4H�4@��#���?                                H�4H�4@                ��+��+@        ��/����?                ��/����?                ��/���@H�4H�4@        ��/����?H�4H�4@                H�4H�4@        ��/����?                ���-��@        ��#�� @                        ��/���@�C=�C=<@                #0#06@        ��/���@H�4H�4@        ��/����?H�4H�4@        ��/����?0#0# @                0#0# @        ��/����?                        0#0#@        �cp>@        ��#��@                z�5��@���-��@�;�;K@        0����/@��8��8J@        0����/@0#0#0@        ��/���@0#0# @        ��/���@0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                �cp>@                        0#0#�?        ��/����?�C=�C=,@        ��/����?�C=�C=@        ��/����?                        �C=�C=@                �C=�C=@                vb'vb'B@                H�4H�4@                B�A�@@z�5��@��/����?0#0# @z�5��@��/����?                ��/����?        z�5��@                                0#0# @�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJUehFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK煔h��B�2         �                  b?�b��S�?/      |�]z}@       �                 ��1�?����tY�?�       ����%)w@       �                  e�?l[jL�?�       ���a�Yq@                          ҏ�?r�8���?�       *���p@                        @���?rF�F!�?       󃥰�G@                        pG�l?�FS�5�?       ��9ՇB@                         h��?4=�%�?       t=�x�-@������������������������       �               ���-��@	                        � Q?����?       ��X�)B @
                        ;��?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?                        P��?      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@                        PP�?��k���?       D+զm76@������������������������       �      ��
       D�JԮD1@                        0�~�?4=�%�?       �(J��@������������������������       �               ��#�� @������������������������       �               �cp>@                         p��?0A����?       4E���_"@                        0��?\����?       P	K��@������������������������       �               ��/����?������������������������       �               z�5��@������������������������       �               0#0# @       S                 �Pv�?��e���?�       *�h�Lvk@       R                 0=T�?*�]����?I       �,^��[@       A                  �E�?�3jG�?B       XC1[+�X@       @                 �j"�?H����?/       ����e�Q@       ;                 �C>?0�<���?.       ��r�MxQ@                         �<��>5�7V��?%       z� �M@������������������������       �               �cp>@!       8                 �!�?B�4w��?$       
��^L@"       5                 �U�?V�%�,�?!       ˠ�I�J@#       4                 �m?l\Cl[��?       @�s�d�I@$       /                  ��~�?����H�?       5���A@%       *                 `q��?P�s�	�?       f���:@&       )                 ��Hb?0 ����?       0
C>�5@'       (                 �_?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �      ��	       ��#��0@+       ,                 �F܂?�d�$���?       �T�f@������������������������       �               ��#�� @-       .                 ��li?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?0       1                  ���?� �_rK�?       J�@��"@������������������������       �               �cp>@2       3                ����t?�����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?������������������������       �        	       �P^Cy/@6       7                 ��2�?j�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?9       :                 ���?~%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?<       =                 D�`?���I@�?	       �2d�%@������������������������       �      ��       �cp>@>       ?                 ��Cw?ܗZ�	7�?       j~���@������������������������       �               z�5��@������������������������       �      �<       ��/����?������������������������       �     ��<       0#0# @B       K                 �]t?�������?       �v���;@C       H                   +Y�?\n����?       Ӏh��K.@D       E                 X[cp?0�c3���?       �uk��!@������������������������       �               ��/���@F       G                 x^��?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?I       J                  �Mm�?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ;��,��@L       Q                 ����?�����?       �l�C�J)@M       N                  �^��?�^�#΀�?       O�{��A%@������������������������       �               ���-��@O       P                 �b'�?��fm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               \Lg1��&@T       {                  ����?��FJ)��?D       k�s��'[@U       d                 �m��?��`$��?.       yn��*R@V       [                 ��@�?1���S��?       KC�S�>@W       Z                 ��aӾ����?       �Ä�>c(@X       Y                 �?
4=�%�?       �(J��@������������������������       �               ��#�� @������������������������       �               �cp>@������������������������       �      ��       ���>��@\       _                  �Q�?��G�%�?       \��rs2@]       ^                 �m۶?z�G���?       '5L�`�@������������������������       �               �cp>@������������������������       �               H�4H�4@`       a                 p:��?��c`�?       %��t5)@������������������������       �      ��       鰑%@b       c                    �?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?e       x                 @��?>�b�% �?       L��_��D@f       s                  @mj�?�uE�~q�?       �ʷ��B@g       p                 P
�?��7m�?       �(�+4@h       o                  _E?`����?       $c�Z%K1@i       n                    �?M�����?       p����.@j       m                 p`�?���/��?       V��7�@k       l                 h�Ѳ?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      �<       ��/����?������������������������       �      ��       [Lg1��&@������������������������       �      ȼ       ��/����?q       r                �I�s?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?t       u                 (�?�p�o䳻?
        9�F�1@������������������������       �               ��#�� @v       w                  ��?�wV����?       Bi�i�"@������������������������       �               0#0#�?������������������������       �               ��#�� @y       z                 p웟?�fm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@|       }                   ���?>�Vv���?       ��)B@������������������������       �               E�JԮD!@~       �                 pt��?������?       %�h�;@       �                 ����?���eCO�?       y3}�0�5@�       �                 Њ�(?p�^AG��?       �7Ѿ1@�       �                 ���?������?	       ��.�SU-@�       �                 @�C�?�L����?       Yk���>)@������������������������       �               ���-��@�       �                 `#��?\%@�"�?       ��[�@������������������������       �               ��#�� @������������������������       �      ��       ��/���@�       �                  ���?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?�       �                 ��j?^����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?�       �                 ����?      �<       ��/���@������������������������       �               ��/����?������������������������       �               �cp>@�       �                 ����?�D#���?       �B�j@������������������������       �               0#0#@������������������������       �               ��#�� @�       �                 ��?Z@G���?	       X��Q'@�       �                 ^7�?z�G���?       '5L�`�@�       �                  P�"�?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �               0#0# @�       �                 \�Z�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               0����/@�       �                   ���?&c4{�"�?9       WM�2�=W@�       �                 ``��?�ݳ��#�?       ��E�b�B@������������������������       �               ;��,��@�       �                 �Q�?
c��rv�?       \����M@@������������������������       �               ���-��@�       �                 P�?w�v1��?        ��O��9@�       �                 pm��? "�7V�?       t	����5@�       �                 X�:�?L� P?)�?       ����x�@������������������������       �               ��#�� @�       �                 ����?T����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @�       �                  �"�?������?       Wؗյ0@������������������������       �               0����/@�       �                 ��	�?��r�g��?       ��1ֻ�'@�       �                  �JV�?�;�a
=�?       ��l��@�       �                   .p�?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?������������������������       �               ��/���@�       �                  Pmj�?L� P?)�?       ����x�@������������������������       �               ��#��@������������������������       �               0#0#�?������������������������       �               0#0#@�       �                  @���?4�>P���?!       �ǒ�a�K@�       �                 �k��?ZJ�ا��?        V�S0f�J@�       �                 @�2�?�J�S��?       ,>���6@�       �                  p�Z?��;�� �?       *.���4@�       �                pnQɠ?�T`�[k�?
       �m����0@�       �                  4�?hutee�?       P9��#@������������������������       �               H�4H�4@������������������������       �      ȼ       ��/���@������������������������       �               �C=�C=@������������������������       �               0#0#@�       �                 `��?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?�       �                 �Y�?d�+(�s�?       ��iq
6>@������������������������       �               ��-��-5@�       �                 ��?�4^��?       s_w$/"@�       �                 �%�?Hy��]0�?       ���y"@������������������������       �               ��/����?������������������������       �               ��+��+@�       �                  `<��?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      �<       ��#�� @�       �                  �E�?ԕFɂ|�?E       �zT��DY@�       �                 @L7�?�L&�ǘ�?%       V�$��I@�       �                 ��Խ?z�G���?
       �'9��1@�       �                 �N��?�� ��?       qp� k'@�       �                 Pn�o?���mf�?       毠�?b#@������������������������       �               0#0# @������������������������       �      �<       ��/���@������������������������       �               0#0# @�       �                  ��d�?Py��]0�?       ���y"@������������������������       �               ��/����?������������������������       �               ��+��+@�       �                 �K�n?����?       bw�ѵA@�       �                 P n?�w��d��?       �0���s@�       �                 Ȑ��?lutee�?       Q9��@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �      �<       ��/����?�       �                 �p�?H�)�n�?       �b�}{.;@������������������������       �      ��       H�4H�48@�       �                 `�m�?���`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 �7T{?H��b�$�?        -�&�H@�       �                 Цt�?�@����?       ���a�#@������������������������       �               0#0# @������������������������       �      ȼ       ��/����?�       �                   ��?      �<       ������C@������������������������       �               �C=�C=@������������������������       �               0#0#@@�t�bh�hhK ��h��R�(KK�KK��h �B�  g:��,&c@�B�)Dd@�dJ�d�c@g:��,&c@����Xb@eJ�dJ�Q@5��t�`@�~Y�u^@��+��+4@5��t�`@G!�M\@S2%S2%1@���>��,@�_��e�=@0#0# @��#�� @��|��<@        z�5��@E�JԮD!@                ���-��@        z�5��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ��#��@                ��#���?                z�5��@                ��#�� @%jW�v%4@                D�JԮD1@        ��#�� @�cp>@        ��#�� @                        �cp>@        z�5��@��/����?0#0# @z�5��@��/����?                ��/����?        z�5��@                                0#0# @r(���F^@[�ڕ��T@�A�A.@�YLg1R@�-����@@��+��+@��>���N@�-����@@��+��+@}�5��H@1����/3@H�4H�4@~�5��H@0����/3@0#0#�?����JG@�cp>'@0#0#�?        �cp>@        ����JG@D�JԮD!@0#0#�?]Lg1��F@���-��@0#0#�?^Lg1��F@�cp>@        Jp�}>@�cp>@        |�5��8@��/����?        <��,��4@��/����?        ��#��@��/����?        ��#��@                        ��/����?        ��#��0@                ��#��@��/����?        ��#�� @                ��#�� @��/����?        ��#�� @                        ��/����?        ;��,��@��/���@                �cp>@        ;��,��@��/����?        ;��,��@                        ��/����?        �P^Cy/@                        ��/����?0#0#�?        ��/����?                        0#0#�?��#���?��/����?                ��/����?        ��#���?                z�5��@��/���@                �cp>@        z�5��@��/����?        z�5��@                        ��/����?                        0#0# @[Lg1��&@��|��,@0#0# @;��,��$@0����/@        ��#��@0����/@                ��/���@        ��#��@��/����?        ��#��@                        ��/����?        z�5��@                ��#���?                ;��,��@                ��#���?0����/#@0#0# @��#���?0����/#@                ���-��@        ��#���?�cp>@                �cp>@        ��#���?                                0#0# @\Lg1��&@                4��tSH@��On�H@��+��+$@=��,��D@���-��:@0#0#@;��,��$@D�JԮD1@H�4H�4@�k(��"@�cp>@        ��#�� @�cp>@        ��#�� @                        �cp>@        ���>��@                ��#���?��|��,@H�4H�4@        �cp>@H�4H�4@        �cp>@                        H�4H�4@��#���?�cp>'@                鰑%@        ��#���?��/����?        ��#���?                        ��/����?        �P^Cy?@/����/#@0#0#�?Jp�}>@���-��@0#0#�?��b:��*@���-��@        ��b:��*@��/���@        ��b:��*@��/����?        ��#�� @��/����?        ��#�� @��/����?        ��#�� @                        ��/����?                ��/����?        [Lg1��&@                        ��/����?                �cp>@                ��/����?                ��/����?        ��#��0@        0#0#�?��#�� @                ��#�� @        0#0#�?                0#0#�?��#�� @                ��#���?�cp>@        ��#���?                        �cp>@        ���>��@�cp>7@H�4H�4@        E�JԮD!@        ���>��@��|��,@H�4H�4@;��,��@��|��,@0#0# @;��,��@鰑%@0#0# @z�5��@鰑%@0#0#�?��#�� @鰑%@                ���-��@        ��#�� @��/���@        ��#�� @                        ��/���@        ��#���?        0#0#�?                0#0#�?��#���?                ��#�� @        0#0#�?��#�� @                                0#0#�?        ��/���@                ��/����?                �cp>@        ��#�� @        0#0#@                0#0#@��#�� @                        D�JԮD!@H�4H�4@        �cp>@H�4H�4@        �cp>@0#0#�?        �cp>@                        0#0#�?                0#0# @        �cp>@                ��/����?                0����/@        ��,���1@��On�8@n�6k�6I@��b:��*@E�JԮD1@�C=�C=@;��,��@                ��#�� @E�JԮD1@�C=�C=@        ���-��@        ��#�� @鰑%@�C=�C=@��#�� @鰑%@H�4H�4@��#��@        0#0#�?��#�� @                ��#�� @        0#0#�?                0#0#�?��#�� @                ��#��@鰑%@0#0# @        0����/@        ��#��@�cp>@0#0# @        �cp>@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/���@        ��#��@        0#0#�?��#��@                                0#0#�?                0#0#@��#��@��/���@�
��
�E@��#�� @��/���@�
��
�E@        �cp>@S2%S2%1@        ��/���@S2%S2%1@        ��/���@��8��8*@        ��/���@H�4H�4@                H�4H�4@        ��/���@                        �C=�C=@                0#0#@        ��/����?                ��/����?                ��/����?        ��#�� @��/����?��8��8:@                ��-��-5@��#�� @��/����?��+��+@        ��/����?��+��+@        ��/����?                        ��+��+@��#�� @��/����?                ��/����?        ��#�� @                ��#�� @                        ��/���.@�~��~nU@        ���-��*@��)��)C@        E�JԮD!@vb'vb'"@        ��/���@0#0#@        ��/���@0#0# @                0#0# @        ��/���@                        0#0# @        ��/����?��+��+@        ��/����?                        ��+��+@        0����/@�s?�s?=@        ��/���@H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@        ��/����?                ��/����?��8��8:@                H�4H�48@        ��/����?0#0# @        ��/����?                        0#0# @        ��/����?7k�6k�G@        ��/����?0#0# @                0#0# @        ��/����?                        ������C@                �C=�C=@                0#0#@@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�)�rhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK߅�h��B�0         ~                 @@�?
��4�?(      ��3�p�}@       ?                   �P�?�*v�o[�?�       I]yQ�9m@       2                 �,�?j]{��`�?N       tF��L^@                        `��?�t�^<{�?A       `ɐ<�6Y@                        �dW?|b8�Y�?       FJͰ(@������������������������       �               ��/����?������������������������       �      �<       [Lg1��&@       )                 �U�<?�5��+'�?<       ���� V@	       (                  �g<�?��U>��?)       m��K��M@
                        ���a?�A&w(�?#       ��|��H@                        ���T?�O-r��?       �.w��e)@                        p�R?�����?       ��X�)B@                        (PH?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?                        0��#?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?������������������������       �               D�JԮD!@                        ��Fo?�.���?       �^���A@������������������������       �               z�5��@       %                 �^Ҧ?6�D��?       �>Dq6/=@       "                 ��r.?�3���r�?       ��7�nN:@                        PRݥ?�d�$���?       �T�f4@                        ౻w?�:V��?       �GP�1@������������������������       �               �k(��"@                        �S�?x�6L�n�?       �E#��h @                        �e?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               z�5��@        !                    �?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?#       $                    �?n%@�"�?       ��[�@������������������������       �      �<       ��/���@������������������������       �               ��#�� @&       '                 �͟�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               �cp>'@*       1                  s��?x�, �#�?       ��
���<@+       .                 �r��?�R�Gz۱?       �P��;@,       -                  ;��?      �<       �cp>�9@������������������������       �               ��/����?������������������������       �               �e�_��7@/       0                 ��u�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      �<       ��#���?3       6                 �mx�?ӝ�h-v�?       N�	��W4@4       5                  ��3�?�_�A�?       肵�e`@������������������������       �               ;��,��@������������������������       �      �<       ��/����?7       >                 ��?�d�����?	       &'9\�~*@8       =                 p۶�?���!��?       �@��&@9       <                ��ߦ�?�D�-,�?       �D'ŰO@:       ;                   E(�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               0#0#@������������������������       �      ȼ       ��/����?������������������������       �               z�5��@@       s                 pL�?��˧��?D       t_�Z&\@A       j                 �@�?p�j�9�?9       {�lW@B       e                 p��?Z�g����?0       ӷ���S@C       \                    �?�uE�~q�?,       �ʷ��R@D       E                 �? M��T��?"       n,��4�N@������������������������       �               ��/����?F       O                 �F��?������?!       �l7�h[N@G       L                  �@r
<`&�?       ���g�F@H       K                 @6�?`�s�	�?       e���*@I       J                 ���>`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               <��,��$@M       N                 `�>      �<       ���b:@@������������������������       �               ��#�� @������������������������       �               Lp�}>@P       Y                 �m.?�K$e_�?	       �EU�}.@Q       T                 ��=�?t����?       ~��qπ*@R       S                  ���?�|2N��?       �3K}@������������������������       �               0#0# @������������������������       �               z�5��@U       X                 �PMT?����?       ��X�)B @V       W                  �G?�?���/��?       V��7�@������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �               ��#��@Z       [                 0p�:?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?]       ^                 �Q�?z�R ��?
       ⲿꁞ+@������������������������       �               ���-��@_       d                ���u?�_�A�?       肵�e`@`       c                  ص�?��Z�	7�?       j~���@a       b                   �x�?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �               ��#�� @f       i                 �>"�?�@G���?       hu��@g       h                 �e�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               0#0#�?k       p                 ��K�?�����?	       Tŵ�)@l       m                 �W�?�֪u�_�?       ��?�8@������������������������       �               �cp>@n       o                 @�g?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?q       r                 ��'�?�.�KQu�?       �K̎@������������������������       �               z�5��@������������������������       �               0#0#@t       u                  ���?���x�?       ��N�H4@������������������������       �               ��+��+@v       y                  �P�?hȃ����?	       1�i?�{.@w       x                 �U�?      �<       ��#�� @������������������������       �               z�5��@������������������������       �               ;��,��@z       {                 `�w?�AP�9��?       i��6��@������������������������       �               H�4H�4@|       }                 hU�<?|�G���?       ��%�|@������������������������       �               0#0# @������������������������       �      �<       ��/����?       �                 ���?�i�	�?�       �:��Y�m@�       �                 p���?,ѝ3� �?C       m��P�k\@�       �                  X?�;f����?'       ?'�'Q@�       �                  ���?I_�+��?       W����<@�       �                 �U��>�~��v��?       ���*@�       �                 �q��?޺W�w��?       �'DQm"@������������������������       �               0#0#�?�       �                 �m�?��6L�n�?       �E#��h @�       �                  ���?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               z�5��@������������������������       �      м       ��/���@�       �                 ���?����|e�?       �z �B�/@�       �                 �U�L?`�ih�<�?       ��
,@�       �                 ��?�n���k�?       3��&�*@�       �                 ��_�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �        	       #0#0&@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?�       �                 0b�?�&��գ�?       PHYCz�C@�       �                 @F�      �<       �C=�C=<@������������������������       �               0#0#�?������������������������       �               �;�;;@�       �                 Pl?�'z�3�?       ���da�%@������������������������       �               H�4H�4@�       �                  2�i?���mf�?       毠�?b@������������������������       �               0#0#�?������������������������       �      �<       ��/���@�       �                 �F�?"�&�Jy�?       X�D}��F@�       �                 T|�?�Ƌ.���?       6U� ��@@�       �                 NK�X?�vL蜇�?       ���>@�       �                 �U�,?rR����?       q\����!@�       �                    �?L� P?)�?       ����x�@������������������������       �               ��#��@������������������������       �               0#0#�?������������������������       �      �<       ��/���@������������������������       �               �k(���5@�       �                 �$�?      �<       H�4H�4@������������������������       �               0#0#�?������������������������       �               0#0# @�       �                 �ڔ?������?       ~���]�'@�       �                 �K�?dQ��?       �s�=�!@������������������������       �      ��       ��/���@�       �                 p���?
4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @������������������������       �               H�4H�4@�       �                 �s�?��0�� �?S       ��NQ�v_@�       �                 ��@s?�����?>       *X�q�X@�       �                 �A�?d�k����?!       �o@ū�F@�       �                 pU�L?R�H�q�?       ��	0�A@�       �                 ���?�w'��h�?       ��,&��4@�       �                 �o�??�?�0�!�?       a`�T�$@������������������������       �               0#0# @�       �                 �Q
�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                    �?&��5�?
       ��~���%@�       �                p�S�?~��j�?       �e��w@�       �                  PV��?T����1�?       ��;9�@������������������������       �               ��#�� @�       �                  ���?�J���?       ��*]Y@������������������������       �               0#0# @������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?������������������������       �      м       ��/���@�       �                 ���?��,���?       !C�s��,@������������������������       �               0����/#@�       �                 ��Z�?���mf�?       毠�?b@������������������������       �               �cp>@�       �                p�K=�?~�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 K��?�?�0�!�?       a`�T�$@������������������������       �               ��/����?������������������������       �               vb'vb'"@�       �                   �?RA���?       �@��J@������������������������       �        
       ��-��-5@�       �                 �Z�?���L�?       >G���@@������������������������       �               ��/����?�       �                   ��?�?�0�!�?       ��G�>@������������������������       �               �C=�C=,@�       �                 �^��?j�q����?       O�Q*s�/@�       �                 0R��?v=���?       � ��R(@������������������������       �               ��/����?������������������������       �               #0#0&@�       �                 ����?v�G���?       ��%�|@������������������������       �               0#0# @������������������������       �      �<       ��/����?�       �                 P��? �)�n�?       �b�}{.;@�       �                 x���?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       k�6k�69@�t�bh�hhK ��h��R�(KK�KK��h �B�  �YLgqd@�-����`@��o���e@�P^Cy_@�H��tXU@H�4H�48@U^CyeJ@2����-O@H�4H�4@��k(/D@�_��e�M@0#0#�?ZLg1��&@��/����?                ��/����?        [Lg1��&@                ���>��<@G�)�BM@0#0#�?,�����;@�]�ڕ�?@        ,�����;@&jW�v%4@        z�5��@0����/#@        z�5��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                ��#���?                ��#���?                        D�JԮD!@        |�5��8@鰑%@        z�5��@                �k(��2@鰑%@        �k(��2@��/���@        ��#��0@��/���@        ��#��0@��/����?        �k(��"@                ���>��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        z�5��@                        �cp>@                ��/����?                ��/����?        ��#�� @��/���@                ��/���@        ��#�� @                        �cp>@                ��/����?                ��/����?                �cp>'@        ��#���?���-��:@0#0#�?        ���-��:@0#0#�?        �cp>�9@                ��/����?                �e�_��7@                ��/����?0#0#�?        ��/����?                        0#0#�?��#���?                z�5��(@�cp>@��+��+@;��,��@��/����?        ;��,��@                        ��/����?        ���>��@��/����?��+��+@��#���?��/����?��+��+@��#���?        ��+��+@��#���?        0#0#�?��#���?                                0#0#�?                0#0#@        ��/����?        z�5��@                ������Q@�cp>7@vb'vb'2@%�}��O@鰑5@0#0# @Lp�}N@On��O0@H�4H�4@Mp�}N@���-��*@0#0# @�>��nK@0����/@0#0# @        ��/����?        �>��nK@��/���@0#0# @�GpAF@��/����?        z�5��(@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        <��,��$@                ���b:@@                ��#�� @                Lp�}>@                <��,��$@�cp>@0#0# @�k(��"@��/����?0#0# @z�5��@        0#0# @                0#0# @z�5��@                z�5��@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ��#��@                ��#���?��/����?                ��/����?        ��#���?                ;��,��@D�JԮD!@                ���-��@        ;��,��@��/����?        z�5��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                ��#�� @                        �cp>@0#0#�?        �cp>@                ��/����?                ��/����?                        0#0#�?z�5��@0����/@��+��+@        0����/@0#0#�?        �cp>@                ��/����?0#0#�?                0#0#�?        ��/����?        z�5��@        0#0#@z�5��@                                0#0#@��#�� @��/����?��+��+$@                ��+��+@��#�� @��/����?��+��+@��#�� @                z�5��@                ;��,��@                        ��/����?��+��+@                H�4H�4@        ��/����?0#0# @                0#0# @        ��/����?        ������C@z%jW�vH@�i��b@��,���A@�cp>7@�+��+�K@���>��@��On�(@H�4H�4H@���>��@D�JԮD!@��8��8*@���>��@0����/@0#0#�?���>��@��/����?0#0#�?                0#0#�?���>��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        z�5��@                        ��/���@                ��/���@H�4H�4(@        ��/����?H�4H�4(@        ��/����?H�4H�4(@        ��/����?0#0#�?        ��/����?                        0#0#�?                #0#0&@        ��/����?                ��/����?                ��/���@dJ�dJ�A@                �C=�C=<@                0#0#�?                �;�;;@        ��/���@�C=�C=@                H�4H�4@        ��/���@0#0#�?                0#0#�?        ��/���@        *�����;@鰑%@�C=�C=@	�#���9@��/���@0#0#@	�#���9@��/���@0#0#�?��#��@��/���@0#0#�?��#��@        0#0#�?��#��@                                0#0#�?        ��/���@        �k(���5@                                H�4H�4@                0#0#�?                0#0# @��#�� @���-��@H�4H�4@��#�� @���-��@                ��/���@        ��#�� @�cp>@                �cp>@        ��#�� @                                H�4H�4@��#��@�cp>�9@B�s?��W@��#��@��On�8@]��[�eQ@��#��@&jW�v%4@��-��-5@��#��@1����/3@H�4H�4(@��#��@�cp>@#0#0&@        ��/����?vb'vb'"@                0#0# @        ��/����?0#0#�?        ��/����?                        0#0#�?��#��@0����/@0#0# @��#��@��/����?0#0# @��#��@        0#0# @��#�� @                ��#�� @        0#0# @                0#0# @��#�� @                        ��/����?                ��/���@                ���-��*@0#0#�?        0����/#@                ��/���@0#0#�?        �cp>@                ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?vb'vb'"@        ��/����?                        vb'vb'"@        0����/@I�4H�4H@                ��-��-5@        0����/@�;�;;@        ��/����?                �cp>@�;�;;@                �C=�C=,@        �cp>@��8��8*@        ��/����?#0#0&@        ��/����?                        #0#0&@        ��/����?0#0# @                0#0# @        ��/����?                ��/����?��8��8:@        ��/����?0#0#�?        ��/����?                        0#0#�?                k�6k�69@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJX"4qhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKӅ�h��B(.         �                 ����? ���7�?%      \4��9{}@       3                 ��Bt?��eJr��?       k�6j/iz@       "                 `%�7?./�o���?F       ��#�O_@                         �\�?�h���a�?3       -���V@                        ~`���:<��?       +:M_Z�4@������������������������       �               0����/#@       
                  `�J�?����X��?       &��֞&@       	                  �q�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       �k(��"@                         ���?xs��?&       ~��`+�Q@                        `f��>�q�Ptܳ?       T�� 5�G@                        ���?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@                        8Q�S?�V_�"�?        ����E@                        P�_?`n����?       � ��w<@������������������������       �               ��#���?                        �U�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?                          ��?      �<       ��k(/D@������������������������       �               ;��,��@������������������������       �               ��,���A@                        x5W�? Xb���?       N�EBCZ7@                        �y������cE��?
       b�co5@                        ؿk?d%@�"�?       ��[�@������������������������       �      ��       ��/���@������������������������       �               ��#�� @������������������������       �      ��       �P^Cy/@        !                 �=��?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?#       *                 �<�?��߭Q��?       �QVl�@@$       %                 ��]?�ۜ�x�?       d��إV3@������������������������       �               E�JԮD!@&       '                 �S�?V�ђ���?       �oFݜh%@������������������������       �               E�JԮD!@(       )                ��f>Y?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?+       .                 ��^?�_�A�?       炵�e`,@,       -                 l�Wr?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?/       0                  p�:?��t� �?       ����x&@������������������������       �               ��/����?1       2                 �@~b?�FO���?       �ߌ$@������������������������       �      ��       �k(��"@������������������������       �      ȼ       ��/����?4       �                 ��?h�xq��?�       .6;aA�r@5       >                  �!�?D�۹C�?�       :3e.6Jl@6       9                   B�?v�����?       u����&:@7       8                 ��?�� N��?
       �L�EBC3@������������������������       �        	       :l��F:2@������������������������       �      �<       ��#���?:       =                  �{��?n��w��?       ���@;       <                 dѬ�?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?������������������������       �               ��/���@?       �                 �6j}?ïBj]��?z       	��tVi@@       �                 �҆�?'�C���?e       �nCe@A       z                 ��&�?��g���?]       ��z���c@B       a                 �A(�?{d�$�?N       ���r_@C       J                 ����?.��V��?)       ����,O@D       I                 <���?�d�$���?       �T�f$@E       F                 ]E?X�j���?       ���z"@������������������������       �               z�5��@G       H                 ��Q?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?K       V                   �x�?���d��?"       �
/�oJ@L       S                 \F�M?   ���?       ,x�1�9@M       N                 �%s?L�r{��?
       e�6� /@������������������������       �               ��#���?O       R                 P�Y�?��&���?	       ��G2��,@P       Q                 ���v?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               �cp>'@T       U                  �~��?      �<       ;��,��$@������������������������       �               ��#���?������������������������       �               �k(��"@W       `                 ��|�?xe�|�/�?       ���f�L:@X       Y                 n�
Q?�����?       �l�C�J9@������������������������       �               ��/���.@Z       _                 p�~�?��`i��?       �؛.�#@[       \                 ��*r?�3`���?       .�r�� @������������������������       �               0#0#@]       ^                   ���?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?������������������������       �               0#0#�?b       o                  ��?�Ojմ��?%       �_���O@c       f                  ��?�4O��?       ���]��9@d       e                 ػ�?�ctn�0�?       �$�k�K @������������������������       �               z�5��@������������������������       �      ��       ��+��+@g       j                 �?�?��íxq�?       �%�'��1@h       i                  ��g�? ܜ�x�?       d��إV#@������������������������       �               E�JԮD!@������������������������       �      �<       ��#���?k       l                 �]�?�̥Q)�?       �9C�<�@������������������������       �               ��#�� @m       n                 `U�?z�G���?       '5L�`�@������������������������       �               H�4H�4@������������������������       �               �cp>@p       u                 uP�?�ti9��?       ��>��B@q       r                 0�~�?�oH2.w�?       �їD́%@������������������������       �               0#0#�?s       t                  ��?& k�Lj�?       �q��l}#@������������������������       �               ��#�� @������������������������       �               ��/���@v       w                 0?���D`|�?       -&ۿ�:@������������������������       �      ��	       �P^Cy/@x       y                 h�B?l7Y���?       ���r�&@������������������������       �               0#0#�?������������������������       �               <��,��$@{       ~                 P�!z?��r�S�?       �f��%?@|       }                   �G�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@       �                  կ?���C��?       >W=��;@������������������������       �               ��|��,@�       �                 0I��?�m:�4�?       ���-X)@������������������������       �               0����/#@�       �                    �?T����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @�       �                 @���?T[�Jg�?       X�S0f�*@������������������������       �               �k(��"@�       �                  ���?E��NV=�?       �t�ܲ@�       �                 ����?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                  ��^�?��E�B��?       eߞKC>@������������������������       �        
       0#0#0@�       �                 @��?�AP�9��?       i��6��+@������������������������       �               vb'vb'"@�       �                  �G?�?���mf�?       寠�?b@������������������������       �      ��       ��/���@������������������������       �               0#0#�?�       �                 �U��?��mG~��?3       dr"(��Q@�       �                 ��\�?����:�?&       ���%�wI@�       �                 �Ys�?���rc�?       �LK���<@�       �                  �"�?���@��?       �<��9@������������������������       �               ��/����?�       �                 �8Ul? v=���?       � ��R8@�       �                 (Y��?��H�&p�?	       L^�3��%@�       �                 �\�?�?�0�!�?       a`�T�$@������������������������       �               vb'vb'"@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?������������������������       �        	       ��8��8*@�       �                 0�!�?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@�       �                 `}��?D�&�=�?       =d���5@�       �                 �6SZ?Y���a�?       �z���2@�       �                 0�q�?>�Z���?       \֎V��-@�       �                  �JV�?��n��?       �-H�\@�       �                 0K�?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �      ��       0����/@�       �                 �?��?>9�)\e�?       `���b @�       �                  @��?      �<       ;��,��@������������������������       �               ��#���?������������������������       �               ��#��@������������������������       �               �cp>@�       �                 ��>�?����|e�?       �z �B�@�       �                  �^��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               0#0# @������������������������       �      ȼ       z�5��@�       �                 `��?�?�0�!�?       a`�T�4@������������������������       �               ��/����?�       �                  ��?8L�0�h�?       k�e�3@������������������������       �      ��
       �A�A.@�       �                 �V�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                 ����?�5��Ɉ�?%       ��#R�H@�       �                 �m�?�^�F�M�?       ~'�5�@@�       �                 0\?�Jn�� �?       �+�i�0@�       �                 ����?|��`p��?       f;3@��!@������������������������       �               0#0#@�       �                 PR��?l�4���?       �tCP��@������������������������       �               �cp>@������������������������       �               0#0# @������������������������       �               0#0# @�       �                  �!�?      �<       0#0#0@������������������������       �               0#0#�?������������������������       �        
       �A�A.@�       �                 ��?L�4X��?       �<�?p�/@�       �                �T�?D��NV=�?       �t�ܲ@�       �                 ��˜?d%@�"�?       ��[�@������������������������       �               ��#���?�       �                 ����?$ k�Lj�?       �q��l}@�       �                 `h�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               0#0# @������������������������       �               0#0# @�t�b�4"     h�hhK ��h��R�(KK�KK��h �B�  u�}e@鰑e@J`F`�`@Qg1���d@��B�)Dd@2��-�rW@����bzU@������C@        ��Gp_R@;l��F:2@        <��,��$@鰑%@                0����/#@        <��,��$@��/����?        ��#���?��/����?                ��/����?        ��#���?                �k(��"@                $�}��O@��/���@        ^Lg1��F@��/����?        z�5��@��/����?                ��/����?        z�5��@                ���#8E@��/����?        ��#�� @��/����?        ��#���?                ��#���?��/����?        ��#���?                        ��/����?        ��k(/D@                ;��,��@                ��,���A@                ��,���1@�cp>@        ��,���1@��/���@        ��#�� @��/���@                ��/���@        ��#�� @                �P^Cy/@                        ��/����?                ��/����?                ��/����?        z�5��(@鰑5@        ��#�� @D�JԮD1@                E�JԮD!@        ��#�� @D�JԮD!@                E�JԮD!@        ��#�� @                ��#���?                ��#���?                <��,��$@��/���@        ��#���?��/����?        ��#���?                        ��/����?        �k(��"@��/����?                ��/����?        �k(��"@��/����?        �k(��"@                        ��/����?        ��k(/T@��/���^@5��-�rW@������Q@��18�Z@H�4H�4H@��#�� @h
��6@0#0# @��#���?:l��F:2@                :l��F:2@        ��#���?                ��#���?��/���@0#0# @��#���?        0#0# @                0#0# @��#���?                        ��/���@        j1��tVQ@鰑U@(S2%S2G@j1��tVQ@'jW�v%T@��+��+4@    �M@������S@��)��)3@u�}wL@���-��J@�A�A.@\Lg1��6@F�JԮDA@��+��+@��#�� @��/����?        ��#�� @��/����?        z�5��@                ��#�� @��/����?                ��/����?        ��#�� @                        ��/����?        ���>��,@On��O@@��+��+@{�5��(@���-��*@        ��#�� @���-��*@        ��#���?                ��#���?���-��*@        ��#���?��/����?        ��#���?                        ��/����?                �cp>'@        ;��,��$@                ��#���?                �k(��"@                ��#�� @0����/3@��+��+@��#�� @0����/3@0#0#@        ��/���.@        ��#�� @��/���@0#0#@��#�� @��/����?0#0#@                0#0#@��#�� @��/����?                ��/����?        ��#�� @                        ��/����?                        0#0#�?Ey�5A@0����/3@��+��+$@z�5��@�cp>'@0#0# @z�5��@        ��+��+@z�5��@                                ��+��+@z�5��@�cp>'@H�4H�4@��#���?D�JԮD!@                E�JԮD!@        ��#���?                ��#�� @�cp>@H�4H�4@��#�� @                        �cp>@H�4H�4@                H�4H�4@        �cp>@        *�����;@��/���@0#0# @��#�� @��/���@0#0#�?                0#0#�?��#�� @��/���@        ��#�� @                        ��/���@        �#���9@        0#0#�?�P^Cy/@                <��,��$@        0#0#�?                0#0#�?<��,��$@                ��#�� @��On�8@0#0#@        ��/����?H�4H�4@        ��/����?                        H�4H�4@��#�� @�e�_��7@0#0#�?        ��|��,@        ��#�� @0����/#@0#0#�?        0����/#@        ��#�� @        0#0#�?                0#0#�?��#�� @                ;��,��$@��/����?0#0#�?�k(��"@                ��#���?��/����?0#0#�?��#���?        0#0#�?                0#0#�?��#���?                        ��/����?                ��/���@��8��8:@                0#0#0@        ��/���@��+��+$@                vb'vb'"@        ��/���@0#0#�?        ��/���@                        0#0#�?�k(��"@Nn��O0@;�;�F@�k(��"@��|��,@�;�;;@        �cp>@%S2%S27@        �cp>@#0#06@        ��/����?                ��/����?#0#06@        ��/����?vb'vb'"@        ��/����?vb'vb'"@                vb'vb'"@        ��/����?                ��/����?                        ��8��8*@        �cp>@0#0#�?                0#0#�?        �cp>@        �k(��"@D�JԮD!@0#0#@z�5��@E�JԮD!@0#0#@z�5��@��/���@0#0#�?��#���?0����/@0#0#�?��#���?        0#0#�?                0#0#�?��#���?                        0����/@        ;��,��@�cp>@        ;��,��@                ��#���?                ��#��@                        �cp>@                ��/����?H�4H�4@        ��/����?0#0#�?        ��/����?                        0#0#�?                0#0# @z�5��@                        ��/����?vb'vb'2@        ��/����?                ��/����?vb'vb'2@                �A�A.@        ��/����?H�4H�4@        ��/����?                        H�4H�4@��#�� @���-��@��+��+D@        �cp>@�A�A>@        �cp>@�C=�C=,@        �cp>@H�4H�4@                0#0#@        �cp>@0#0# @        �cp>@                        0#0# @                0#0# @                0#0#0@                0#0#�?                �A�A.@��#�� @��/���@��+��+$@��#�� @��/���@0#0# @��#�� @��/���@        ��#���?                ��#���?��/���@        ��#���?��/����?                ��/����?        ��#���?                        �cp>@                        0#0# @                0#0# @�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ;�3whFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK煔h��B�2         �                 ��\�?&]IcQ�?-      ��A=��}@       �                 n~?�n6�$�?�       ���b�q@       p                 P�}A?���W�?�       ����)p@       o                 �J��?�����?z       ��v��h@       &                 X\ ?d��=��?y       �����Zh@                         ��m?4a(���?'       3��h��L@                        �7�<?�'����?       W��Fx�:@                          ���?p%@�"�?       Ͱrɱ�-@	       
                 `���>p@ȱ��?	       pm���S'@������������������������       �               ��#���?                          ��?�^�#΀�?       N�{��A%@������������������������       �      ��       ���-��@                        :�1�>Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?                       @S.�#?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ��#�� @                        0M>c?�����?       �Ä�>c(@                         P�J�?��t� �?       ����x&@                        �r��?�FO���?       �ߌ$@������������������������       �               �k(��"@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?������������������������       �      м       ��/����?       %                 P��1?�FO���?       ,��N�>@       "                    �?|�6L�n�?       ��4}i�8@                        ���}?�hK)�?       �h��K�2@������������������������       �      ��       <��,��$@       !                 �
Y?��6L�n�?       �E#��h @                         ��?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      �<       ;��,��@#       $                  ����?Zn����?       � ��w<@������������������������       �               ��#��@������������������������       �      �<       ��/����?������������������������       �               z�5��@'       B                 P�p�?�2��ˍ�?R       -��!a@(       9                 ��yh?ycP�Fc�?       D��[߲H@)       6                 p۶�?VJ����?       
�CC�<@*       +                 ��5P?��o��^�?       NjO���5@������������������������       �               ;��,��@,       5                 .25Q?ʳI3�?       ���0@-       0                  E(�?D
:����?       |��"�%@.       /                 p��h?�����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?1       2                 �vq?���mf�?       毠�?b@������������������������       �               ��/����?3       4                 �J�{?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �      ��       �cp>@7       8                 �py?d�ih�<�?       ��
@������������������������       �               ��/����?������������������������       �               H�4H�4@:       =                      �3��F��?       nf9t{y4@;       <                 p�լ?      �<
       ��#��0@������������������������       �               ��#���?������������������������       �        	       �P^Cy/@>       A                  ����?̔fm���?       ��Z�N@?       @                 �j%?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��#���?C       N                 ��=�?Z�* �\�?3       <�%��U@D       E                 @+{�?� �^�?�?       ���[r9@������������������������       �               ��On�(@F       M                �E9�?��z}-�?       ��(�I�)@G       J                 �Ι?�*P��?       �����&@H       I                  Џ~�?�����?       ��X�)B @������������������������       �               ��/����?������������������������       �      �<       z�5��@K       L                  н��?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?������������������������       �      м       ��/����?O       T                 �=��?�����?&       �<�OfO@P       Q                   ���?�FO���?       �ߌ$@������������������������       �      ��       ��#�� @R       S                 �!�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?U       V                  bx�?^fG��?        ��/�.�I@������������������������       �               0����/@W       l                 P
�?^P�]��?       /�Ϸ2�G@X       Y                 �j��?�3���r�?       W�i�ҺC@������������������������       �               ��/���@Z       a                    �?nU�vѢ�?       lӶ��A@[       \                 0��?Hn����?       ~��Y-2@������������������������       �               �cp>@]       `                  �g<�?�d�$���?
       ;��#�.@^       _                 �q�3?<9�)\e�?       _���b @������������������������       �               ;��,��@������������������������       �               �cp>@������������������������       �      ȼ       ���>��@b       k                 ��>?y�<�?       X&b��q1@c       j                 �9�?��t� �?       ����x&@d       g                  `K�?�FO���?       �ߌ$@e       f                �w�(�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @h       i                 З��?      �<       ���>��@������������������������       �               ��#���?������������������������       �               z�5��@������������������������       �      ȼ       ��/����?������������������������       �               z�5��@m       n                �I�s?      �<       ��/���@������������������������       �               �cp>@������������������������       �               0����/@������������������������       �               �cp>@q       t                 �m�?Lʺ�;��?)       ��R��qN@r       s                  p��?����x�?       
�ra6�:@������������������������       �               �cp>�9@������������������������       �               0#0#�?u       �                 pf �?I���Rg�?       愙��@@v       }                 `9�`?t����?	       ��qπ*@w       z                 ȟ�Q?�FO���?       �ߌ$@x       y                  P�"�?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@{       |                 ��=�?      �<       z�5��@������������������������       �               ��#�� @������������������������       �               ��#��@~                        b���?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 ���?`�Jm�?       ��E�ǹ4@�       �                  ���?�F���?	       :�.�-'@������������������������       �               ��#���?������������������������       �      ��       鰑%@�       �                 �J�?���A���?       ��\�F"@�       �                 @���?��b�}�?       ���\�@�       �                 H��?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �               ��#��@�       �                 ��K�?�u=���?       � ��R8@�       �                 h�W�?�AP�9��?       i��6��@������������������������       �               ��+��+@������������������������       �      �<       ��/����?������������������������       �        
       S2%S2%1@�       �                 �-�?o���?|       ��[�,�g@�       �                  ��~�?��h��?K       �9���}[@�       �                 �q�?BG��2�?       ��\]�5@�       �                 ��?ܗZ�	7�?       i~���$@������������������������       �               �cp>@�       �                     �?T����?       P	K��@������������������������       �               ��/����?������������������������       �               z�5��@�       �                   s��?�!�a6Z�?	       ���t0�'@�       �                 �C8�? �Ϟi�?       
��ؠ�!@������������������������       �               0#0#@�       �                   E(�?���mf�?       毠�?b@�       �                 �_��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?�       �                 (-��?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ȼ       �cp>@�       �                 Ш��?����>�?:       }6gZ
V@�       �                 ����?��H�&p�?.       ���Q~P@�       �                   �?�g�\CY�?(       B��(M@�       �                  �E�?�-�bƲ?       >�7*9@�       �                    �?�?�0�!�?	       a`�T�$@������������������������       �               ��+��+@�       �                 ��e�?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?������������������������       �      �<
       �A�A.@�       �                 �ں�?�}�	���?       "�Ռx@@�       �                  �>�?��9 ���?       �z��)�6@�       �                 (d��?h��ճC�?	       y��l$,@������������������������       �               #0#0&@�       �                 �|�?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 �9L�?�� ��?       U?
@�!@������������������������       �               �cp>@������������������������       �               H�4H�4@������������������������       �               ��+��+$@�       �                  `���?��G���?       ��%�|@������������������������       �               0#0# @�       �                 P�l�?�� ��?       qp� k@������������������������       �               �cp>@�       �                 AW�?x��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 �@�?      �<       #0#06@������������������������       �               0#0# @������������������������       �               ��+��+4@�       �                 ����?2����?1       �;*�g�S@�       �                 ��?^���f"�?*       >äD�RQ@�       �                 �ܣe?X3��j��?%       	_h�(N@�       �                 `�C?��!�	m�?       A�^�%G@�       �                 pb)�?�[����?       ,�"�o�A@�       �                 ��? �k����?       b*pn�4@�       �                 @�[�?��h��?       S�D'�@������������������������       �               ��#��@�       �                 Ȉ.�?�D#���?       �B�j@������������������������       �               0#0#�?�       �                 03��?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               ��b:��*@�       �                 ����?@o��IF�?       ����	.@�       �                 _%?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0# @������������������������       �               ���>��@�       �                 @� �?�^�#΀�?       O�{��A%@�       �                    �?      �<       /����/#@������������������������       �               ��/���@������������������������       �               �cp>@������������������������       �      ܼ       ��#���?�       �                 ��M�?��ih�<�?	       ��
,@�       �                  ��?lutee�?       Q9��@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               vb'vb'"@�       �                   ���?d����?       �����!@�       �                 P�$�?|�G���?       ��%�|@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �      ��       ��+��+@�       �                 ���?      �<       ��+��+$@������������������������       �               0#0#�?������������������������       �               vb'vb'"@�t�bh�hhK ��h��R�(KK�KK��h �B�  �YLgqd@c
���c@�z��z�b@�P^CyM`@�����]@T2%S2%A@�P^CyM`@�@S4]@H�4H�4(@v�}w\@t�'�x�R@0#0# @v�}w\@=l��F:R@0#0# @���#8E@��/���.@        ���>��,@��On�(@        ;��,��@/����/#@        ��#�� @0����/#@        ��#���?                ��#���?/����/#@                ���-��@        ��#���?�cp>@                �cp>@        ��#���?                z�5��@                ��#���?                ��#�� @                �k(��"@�cp>@        �k(��"@��/����?        �k(��"@��/����?        �k(��"@                        ��/����?                ��/����?                ��/����?        ,�����;@�cp>@        �k(���5@�cp>@        ��,���1@��/����?        <��,��$@                ���>��@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ;��,��@                ��#��@��/����?        ��#��@                        ��/����?        z�5��@                ������Q@��|��L@0#0# @+�����;@��|��,@�C=�C=@;��,��$@�cp>'@�C=�C=@<��,��$@鰑%@0#0#�?;��,��@                ;��,��@鰑%@0#0#�?;��,��@0����/@0#0#�?;��,��@��/����?        ;��,��@                        ��/����?                ��/���@0#0#�?        ��/����?                ��/����?0#0#�?                0#0#�?        ��/����?                �cp>@                ��/����?H�4H�4@        ��/����?                        H�4H�4@��,���1@�cp>@        ��#��0@                ��#���?                �P^Cy/@                ��#���?�cp>@                �cp>@                ��/����?                ��/����?        ��#���?                �k(���E@��]�ڕE@0#0#�?z�5��@:l��F:2@0#0#�?        ��On�(@        z�5��@�cp>@0#0#�?z�5��@��/���@0#0#�?z�5��@��/����?                ��/����?        z�5��@                        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?        �k(��B@��On�8@        �k(��"@��/����?        ��#�� @                ��#���?��/����?        ��#���?                        ��/����?        ,�����;@�e�_��7@                0����/@        ,�����;@0����/3@        ,�����;@�cp>'@                ��/���@        ,�����;@��/���@        z�5��(@�cp>@                �cp>@        {�5��(@�cp>@        ;��,��@�cp>@        ;��,��@                        �cp>@        ���>��@                �P^Cy/@��/����?        �k(��"@��/����?        �k(��"@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ���>��@                ��#���?                z�5��@                        ��/����?        z�5��@                        ��/���@                �cp>@                0����/@                �cp>@        ��#��0@&jW�v%D@0#0#@        �cp>�9@0#0#�?        �cp>�9@                        0#0#�?��#��0@��|��,@H�4H�4@�k(��"@��/����?0#0# @�k(��"@��/����?        z�5��@��/����?                ��/����?        z�5��@                z�5��@                ��#�� @                ��#��@                        ��/����?0#0# @        ��/����?                        0#0# @���>��@��On�(@0#0#�?��#���?鰑%@        ��#���?                        鰑%@        z�5��@��/����?0#0#�?��#�� @��/����?0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?        ��#�� @                ��#��@                        ��/����?#0#06@        ��/����?��+��+@                ��+��+@        ��/����?                        S2%S2%1@��#��@@�)�B�D@�[��[�\@z�5��@h
��6@�N��NlT@z�5��@鰑%@��+��+@z�5��@��/���@                �cp>@        z�5��@��/����?                ��/����?        z�5��@                        ���-��@��+��+@        ��/���@��+��+@                0#0#@        ��/���@0#0#�?        �cp>@                ��/����?                ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@                �cp>'@��)��)S@        �cp>'@�;�;K@        ��/���@j�6k�6I@        ��/����?H�4H�48@        ��/����?vb'vb'"@                ��+��+@        ��/����?0#0#@                0#0#@        ��/����?                        �A�A.@        ���-��@��8��8:@        ���-��@0#0#0@        ��/����?��8��8*@                #0#0&@        ��/����?0#0# @        ��/����?                        0#0# @        �cp>@H�4H�4@        �cp>@                        H�4H�4@                ��+��+$@        ��/���@0#0#@                0#0# @        ��/���@0#0# @        �cp>@                ��/����?0#0# @        ��/����?                        0#0# @                #0#06@                0#0# @                ��+��+4@��b:��:@/����/3@B�A�@@��b:��:@/����/3@%S2%S27@��b:��:@D�JԮD1@0#0#0@��b:��:@��/���.@0#0#@�#���9@�cp>@0#0#@�k(��2@        0#0# @;��,��@        0#0# @��#��@                ��#���?        0#0# @                0#0#�?��#���?        0#0#�?��#���?                                0#0#�?��b:��*@                ���>��@�cp>@0#0# @        �cp>@0#0# @        �cp>@                        0#0# @���>��@                ��#���?/����/#@                /����/#@                ��/���@                �cp>@        ��#���?                        ��/����?H�4H�4(@        ��/����?H�4H�4@        ��/����?                        H�4H�4@                vb'vb'"@        ��/����?�C=�C=@        ��/����?0#0# @                0#0# @        ��/����?                        ��+��+@                ��+��+$@                0#0#�?                vb'vb'"@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�3hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK텔h��B�3         �                  t0�?��I�P�?%      7�	�x}@       �                  ���?z:��uV�?�       a��,ߐu@       :                 pb��?n�>���?�       �-��yq@       3                 �eU�?‥�)R�?U       �1�Ma@       (                 �:W>?N.�L�?N        }I�`@       '                 p5W�?�3,���?;       �r���X@                           �?�qr�Ml�?:       �Se��W@       	                  �Ԧ�?������?&       ���ѫO@������������������������       �               �cp>@
                        �Ԏ?���`�^�?$       +Z�6m;N@                        `�լ?C	���?       �$r.X{?@                         ����?����X��?       '��֞&@������������������������       �               ��/����?������������������������       �      �<       <��,��$@                        ,*�����7m�?
       �(�+4@                         �3��?Ȕfm���?       ��Z�N@������������������������       �               ��#�� @������������������������       �               �cp>@                        x��?|b8�Y�?       FJͰ(@������������������������       �               ��/����?������������������������       �               [Lg1��&@������������������������       �               ���>��<@                        �7�<?Zutee�?       ��@@                        @�4�>�`@s'��?       Di_y,*@������������������������       �               ��/���@                        �ޗ?^%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?                          ҏ�?nzw��?       �B޳�X9@������������������������       �               �cp>@       $                 ��]"?��t� �?       ����x6@        !                 �p�?� �_rK�?       J�@��"@������������������������       �               z�5��@"       #                 Xy�?d%@�"�?       ��[�@������������������������       �      �<       ��/���@������������������������       �               ��#�� @%       &                 P��p?      �<       ��b:��*@������������������������       �               ��#�� @������������������������       �               ZLg1��&@������������������������       �      �       �cp>@)       0                 p��Y?px�TR�?       ���e>@*       +                  �Q�?4=�%�?       �(J��3@������������������������       �      ��       鰑%@,       /                 �<�?l�j���?       ���z"@-       .                  �_�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      �<       ���>��@1       2                  9��?�}	;	�?       vK�>4%@������������������������       �               0����/#@������������������������       �               0#0#�?4       5                  ���?|ۜ�x�?       d��إV#@������������������������       �      ��       ���-��@6       7                 p�E�?d%@�"�?       ��[�@������������������������       �               ��/����?8       9                  P�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?;       <                 �~�?���m�?V       S\l�`@������������������������       �               0#0#@=       |                 �g��?�ұ��?T       �:�JTj`@>       w                 �m��?�����u�??       MT��.�Y@?       X                 ��>}?
-Y�T�?9       ��>_��W@@       U                  D`�?xH4x J�?       ��e�a�A@A       T                 h��?ߍO����?       �o�h37>@B       Q                 p8L�?Z���=k�?       ��kV;@C       P                 �d?6�y�jR�?       �u�̣u8@D       I                 X��?�n�gn��?       �E��ss7@E       H                 Hq$�?ʔfm���?       ��Z�N@F       G                 P\�>      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��#���?J       M                 ����?�U1��-�?	       8�KY��3@K       L                 h�լ?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @N       O                 ��d?�C=+��?       b��T|0@������������������������       �               ��/����?������������������������       �      ��       �P^Cy/@������������������������       �               0#0#�?R       S                 0���?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �      �<       �cp>@V       W                 pU�<?      �<       �cp>@������������������������       �               ��/���@������������������������       �               ��/����?Y       j                 `y��?�M��ө�?$       ��<��M@Z       e                 �M}C?�skҎA�?       ������B@[       d                 �^5?�(�����?	       ��0��0@\       a                 @8��?p���A�?       2gX\-@]       `                      (��c`�?       %��t5)@^       _                 �ȿ? ܜ�x�?       d��إV#@������������������������       �      ��       D�JԮD!@������������������������       �      �<       ��#���?������������������������       �               �cp>@b       c                  ����?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#�� @f       i                 �ז�?@H�,.̷?
       �J�$r.5@g       h                 p)�? ܜ�x�?       d��إV#@������������������������       �               E�JԮD!@������������������������       �      �<       ��#���?������������������������       �               �cp>'@k       n                 H��?A���}�?       �#��5@l       m                 p�?���mf�?       寠�?b#@������������������������       �      ��       ��/���@������������������������       �               0#0# @o       r                �s�[w? ����?	       �Ä�>c(@p       q                 hU�<?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?s       v                 `&�?X�j���?       ���z"@t       u                    �?      �<       ��#�� @������������������������       �               z�5��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?x       {                 @�X�?�AP�9��?       h��6��@y       z                 @��?Hy��]0�?       ���y"@������������������������       �               ��+��+@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?}       �                 p��I?�\�����?       ���I�<@~       �                 4�?�y���@�?       �+�&�G-@       �                 p۶�?)���?       y��uk!@�       �                 �U��>      �<       ���-��@������������������������       �               ��/���@������������������������       �               �cp>@�       �                  �9��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 pe�?uT �+��?       ��>Y��@�       �                  Pmj�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?�       �                  `���?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@�       �                 @E��?t��ճC�?       y��l$,@�       �                 ~R�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               H�4H�4(@�       �                  a��?�fG
�?+       s+:���Q@�       �                 p���?R������?%       �"�IN@�       �                 p)�J?�����?       l�����G@�       �                 �?e?����?       ���
7@�       �                 `B4b?�FO���?       �ߌ$@������������������������       �               ��#�� @�       �                  �^��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                    �?K�A���?       3����)@�       �                ��O�y?��[����?       Hl�_A@�       �                   B�?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �               0����/@������������������������       �               0#0#�?�       �                 ���?z��`p��?       �����@������������������������       �               ��/����?������������������������       �      ��       0#0#@�       �                 T�Y?      �<       H�4H�48@������������������������       �               0#0#@������������������������       �               ��+��+4@�       �                 p'v�?��w�(�?       Z����*@�       �                    �?�wV����?       Bi�i�"@������������������������       �               z�5��@�       �                  �G?�?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?������������������������       �               0#0#@�       �                 p��?F�ђ���?       �oFݜh%@������������������������       �               ���-��@�       �                 �#�?���/��?       V��7�@������������������������       �      �<       ��/����?������������������������       �               ��#�� @�       �                 h��?8����?O       �7*ǜ_@�       �                 �%��?����9�?1       pVB�:�S@�       �                 �b'�?�5�JvZ�?       ����6�A@�       �                 ���?�N�+�?       ����:@�       �                  �P��?��(v��?	       �A�s(.@�       �                 ��:�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               ��8��8*@�       �                 p��I?���};��?	       ��;̑�%@�       �                 P�d�?x�G���?       '5L�`�@������������������������       �               �cp>@������������������������       �               H�4H�4@������������������������       �               ��+��+@�       �                ���?b%��̫�?       �@�o#@�       �                 �=��?)���?       y��uk!@������������������������       �               ��#���?������������������������       �               ��/���@������������������������       �               0#0#�?�       �                 `Fe�?0ӄ%&�?       @��>F@�       �                 ����?Jy��]0�?       �N-ۙ2@������������������������       �               ��/����?�       �                 �8U|?(r����?
       Qz�i0@�       �                 �/�?|��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �      ��       ��8��8*@�       �                 @X!�?      �<       ��8��8:@������������������������       �               0#0#�?������������������������       �               k�6k�69@�       �                     �?P���.��?       D±�=G@�       �                ����?Hy��]0�?       ���y"@������������������������       �               ��/����?������������������������       �               ��+��+@�       �                  @?��?��'':��?       q�`�<D@�       �                 P�?2k�"O��?       �?<��*&@������������������������       �               z�5��@�       �                 @���?, k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?�       �                 `�3W?,����i�?       ��shd=@�       �                  '
�?�tB���?       hW��v4@�       �                    �?(PThD]�?	       �p�]�*@�       �                 Ш��?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?�       �                  ���?X7Y���?       ���r�&@�       �                  ��?�zœ���?       IG���t@�       �                 @��8?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �               ���>��@������������������������       �               �C=�C=@�       �                 ����?|��`p��?       e;3@��!@�       �                 ����?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �      ��       ��+��+@�t�bh�hhK ��h��R�(KK�KK��h �B8  ���khc@�Y���d@�����b@5��t�`@}����a@<��8�cP@���>��\@`�_���_@�A�A>@�YLgqT@�a#6�K@0#0#�?��k(/T@��h
�G@0#0#�?�YLg1R@�cp>�9@        �YLg1R@�cp>7@        V^CyeJ@鰑%@                �cp>@        T^CyeJ@��/���@        �,����7@��/���@        ;��,��$@��/����?                ��/����?        <��,��$@                ��b:��*@���-��@        ��#�� @�cp>@        ��#�� @                        �cp>@        [Lg1��&@��/����?                ��/����?        [Lg1��&@                ���>��<@                ������3@��On�(@        ��#���?�cp>@                ��/���@        ��#���?��/����?        ��#���?                        ��/����?        �k(��2@���-��@                �cp>@        �k(��2@��/���@        ;��,��@��/���@        z�5��@                ��#�� @��/���@                ��/���@        ��#�� @                ��b:��*@                ��#�� @                ZLg1��&@                        �cp>@        ��#�� @鰑5@0#0#�?��#�� @�cp>'@                鰑%@        ��#�� @��/����?        ��#���?��/����?        ��#���?                        ��/����?        ���>��@                        0����/#@0#0#�?        0����/#@                        0#0#�?��#���?E�JԮD!@                ���-��@        ��#���?��/����?                ��/����?        ��#���?��/����?                ��/����?        ��#���?                Ey�5A@~����Q@�s?�s?=@                0#0#@Ey�5A@}����Q@k�6k�69@���b:@@<��18N@��+��+$@���b:@@F�)�BM@��+��+@��,���1@��/���.@H�4H�4@��,���1@/����/#@H�4H�4@��,���1@���-��@H�4H�4@��,���1@��/���@H�4H�4@��,���1@��/���@0#0# @��#���?�cp>@                �cp>@                ��/����?                ��/����?        ��#���?                ��#��0@��/����?0#0# @��#���?        0#0# @��#���?                                0#0# @�P^Cy/@��/����?                ��/����?        �P^Cy/@                                0#0#�?        �cp>@                ��/����?                ��/����?                �cp>@                �cp>@                ��/���@                ��/����?        ���>��,@��]�ڕE@0#0# @;��,��@On��O@@        ��#��@��On�(@        ��#�� @��On�(@        ��#���?�cp>'@        ��#���?E�JԮD!@                D�JԮD!@        ��#���?                        �cp>@        ��#���?��/����?                ��/����?        ��#���?                ��#�� @                ��#���?&jW�v%4@        ��#���?D�JԮD!@                E�JԮD!@        ��#���?                        �cp>'@        �k(��"@鰑%@0#0# @        ��/���@0#0# @        ��/���@                        0#0# @�k(��"@�cp>@        ��#���?��/����?                ��/����?        ��#���?                ��#�� @��/����?        ��#�� @                z�5��@                ;��,��@                        ��/����?                ��/����?��+��+@        ��/����?��+��+@                ��+��+@        ��/����?                ��/����?        ��#�� @�cp>'@�A�A.@��#�� @鰑%@0#0# @��#���?��/���@                ���-��@                ��/���@                �cp>@        ��#���?��/����?                ��/����?        ��#���?                ��#���?�cp>@0#0# @��#���?        0#0#�?��#���?                                0#0#�?        �cp>@0#0#�?                0#0#�?        �cp>@                ��/����?��8��8*@        ��/����?0#0#�?        ��/����?                        0#0#�?                H�4H�4(@������3@On��O0@eJ�dJ�A@��,���1@��/���@dJ�dJ�A@�k(��"@��/���@�A�A>@�k(��"@��/���@H�4H�4@�k(��"@��/����?        ��#�� @                ��#���?��/����?                ��/����?        ��#���?                        ���-��@H�4H�4@        0����/@0#0# @        0����/@0#0#�?                0#0#�?        0����/@                        0#0#�?        ��/����?0#0#@        ��/����?                        0#0#@                H�4H�48@                0#0#@                ��+��+4@��#�� @        ��+��+@��#�� @        0#0#�?z�5��@                ��#�� @        0#0#�?��#�� @                                0#0#�?                0#0#@��#�� @D�JԮD!@                ���-��@        ��#�� @��/����?                ��/����?        ��#�� @                ������3@h
��6@��-��-U@��#���?��|��,@2#0#P@��#���?�cp>'@%S2%S27@        ��/���@#0#06@        ��/����?�C=�C=,@        ��/����?0#0#�?                0#0#�?        ��/����?                        ��8��8*@        �cp>@0#0# @        �cp>@H�4H�4@        �cp>@                        H�4H�4@                ��+��+@��#���?��/���@0#0#�?��#���?��/���@        ��#���?                        ��/���@                        0#0#�?        �cp>@�ڬ�ڬD@        �cp>@�A�A.@        ��/����?                ��/����?�A�A.@        ��/����?0#0# @                0#0# @        ��/����?                        ��8��8*@                ��8��8:@                0#0#�?                k�6k�69@�k(��2@��/���@��+��+4@        ��/����?��+��+@        ��/����?                        ��+��+@�k(��2@���-��@�A�A.@���>��@��/���@        z�5��@                ��#���?��/���@                ��/���@        ��#���?                [Lg1��&@�cp>@�A�A.@ZLg1��&@        vb'vb'"@[Lg1��&@        0#0# @��#���?        0#0#�?                0#0#�?��#���?                ;��,��$@        0#0#�?z�5��@        0#0#�?��#���?        0#0#�?                0#0#�?��#���?                ��#�� @                ���>��@                                �C=�C=@        �cp>@H�4H�4@        �cp>@0#0#�?                0#0#�?        �cp>@                        ��+��+@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ� �NhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK텔h��B�3         �                 p*��?{��T�P�?.       5'�}@       }                  ���?tiCBГ�?�       �+��oq@       p                 �R�?�,ėW�?�       D:ۻ�+l@       c                 ��x�?�B[d}�?�       �����lj@       >                 ���?�݅����?v       l�]�f@                        ��cn?8�,	%��?Q       ����^@                         nl?`�����?!       镁�3�J@                        �ZS?ΐ��b�?       '}#�D�B@	                         ���?j����?       ;��18>@
                        �ofl?΃�\��?       �D+զm7@                        ���a?��t� �?       ����x6@                        �m۶?h����?
       $c�Z%K1@������������������������       �               �k(��"@                        �c:?���/��?       V��7�@������������������������       �               ��/���@������������������������       �               ��#��@������������������������       �               ;��,��@������������������������       �      �<       ��/����?                        POj"?�`@s'��?       Ei_y,*@������������������������       �               �cp>@������������������������       �               ��#���?                         ��^�?��[����?       Hl�_A@������������������������       �               0����/@������������������������       �               0#0# @                         @?��?�h��%�?
       �1�
�u0@������������������������       �      ��       0����/#@                        0?��|��?       ���ĺw@                        ����?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               �cp>@        =                 ��{�?��ř���?0       �w�|Q@!       0                 (�+0?X�ƈ��?.       ���Q@"       )                 ��u�?��X3��?!       h���I@#       (                 ���p?X���B�?       �(R� A@$       %                  �P��?����?       ��X�)B @������������������������       �               ;��,��@&       '                 �G�o?`%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               �#���9@*       /                 `s5�?�S�l�?
       ��8	+*1@+       ,                 �NZ?���`�?       ��
�Me@������������������������       �               0����/@-       .                 ����?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               �k(��"@1       :                 ��nZ?�A53���?       G����0@2       5                 �|y?ʔfm���?
       �0��z'@3       4                  ��M?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?6       9                  ��?�(���?       y��uk!@7       8                 P.�?f%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �               �cp>@;       <                    �?�|2N��?       �3K}@������������������������       �               z�5��@������������������������       �               0#0# @������������������������       �      �       ��/����??       P                 �6F�?��d]P�?%       �+�V��J@@       M                    �?j�n3��?       ś2��4@A       L                  ���?Zn����?       Ӏh��K.@B       G                 ���b?���/��?       5��o��#@C       D                 �/��?�d�$���?       �T�f@������������������������       �               ��/����?E       F                 �)�H?      �<       ��#��@������������������������       �               ��#�� @������������������������       �               ��#�� @H       I                 ��Ɲ?  k�Lj�?       �q��l}@������������������������       �               �cp>@J       K                 ��Lr?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ��       ;��,��@N       O                  ��d�?t@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@Q       Z                 ��܌?f���b��?       �ݧ]@$@@R       S                 �p��?����X�?       ��\M7@������������������������       �               ���-��*@T       W                 0���?XV�IS��?       (���d�#@U       V                �J��?��Z�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@X       Y                  "��?���mf�?       毠�?b@������������������������       �      �<       ��/���@������������������������       �               0#0#�?[       \                 ��-�?��Zu��?       �%���!@������������������������       �               ��/����?]       b                 ����?��G9�?       ���=A@^       _                 �UaG?�@����?       ���a�@������������������������       �               H�4H�4@`       a                 �,��?x�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               ��#�� @d       e                 ��r<?�ޝ  ~�?       P@��WA@������������������������       �               ��/����?f       o                 ���?l��e��?       [��%b@@g       n                    �?�L�����?       p����>@h       m                   �0�?�3���r�?       ��7�nN*@i       l                 PeT�?��t� �?       ����x&@j       k                 `U�?��Z�	7�?       j~���@������������������������       �               z�5��@������������������������       �      �<       ��/����?������������������������       �      ��       z�5��@������������������������       �      ȼ       ��/����?������������������������       �               ��,���1@������������������������       �               0#0# @q       |                 �6Jy?���1p8�?	       |곯�+@r       w                 � K�?f�B��#�?       I[���%@s       v                 ����?��íxq�?       %2��-�@t       u                  н��?���mf�?       寠�?b@������������������������       �      ��       ��/���@������������������������       �               0#0#�?������������������������       �               ��#���?x       y                   �P�?�o���?       o�9�F@������������������������       �               0#0# @z       {                 �ʨ�?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?������������������������       �               H�4H�4@~       �                 ���U?�~*)��?!       bs9��J@       �                 ���>��oR��?       m�Q6�(@������������������������       �               ��/����?�       �                 0�Έ?l7Y���?       ���r�&@������������������������       �               �k(��"@�       �                    �?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?�       �                  �^�?��͈-��?       9��$�D@�       �                 @�V�?O6��j�?       ?Sv�1@�       �                 ��?�C>�?       �1�m�!@������������������������       �               �cp>@�       �                  p�?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?�       �                 ��5�?x�t1u�?       "�te!� @������������������������       �      ��       ���>��@������������������������       �               0#0#�?�       �                 0��?��ߜ���?       �2Ӂ58@�       �                 ��u�?H,�#6?�?       ���*4@�       �                 n�
Q?�v�;B��?       ՟���	 @������������������������       �               ��/����?������������������������       �               �C=�C=@������������������������       �      ��       H�4H�4(@�       �                 ���?�J���?       ��*]Y@������������������������       �               0#0# @������������������������       �               ��#�� @�       �                 ��?�50g�?y       8.�}"h@�       �                 л��?Hk/����?F       r�w[@�       �                  �~��?�ና���?3       q7���S@�       �                 ����?\^�R1�?       H;9X@@�       �                 аs}?fd_Јn�?       ,4���2@�       �                 ��#�?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @�       �                 �vs�?����w�?
       ���Ã@/@�       �                  ��?& k�Lj�?	       d*�}#<-@�       �                 @? ��c`�?       %��t5)@�       �                  'V�?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               /����/#@������������������������       �               ��#�� @������������������������       �               0#0#�?������������������������       �      �<
       ��|��,@�       �                 ����?<�0u��?       �3w�?�F@�       �                 @��?:Y�c�?       �e7#J�=@������������������������       �               H�4H�4@�       �                 �2*�?~i�O��?       U�0���:@�       �                 @�C�?�� �6�?	       ���*9�0@�       �                 ��ɬ?��^���?       ���w!@�       �                 p���?d�4���?       �tCP��@�       �                   +Y�?���`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               ��/���@�       �                 0.��?@9�)\e�?       _���b @������������������������       �               ;��,��@������������������������       �               �cp>@�       �                  ��d�?jutee�?       Q9��#@������������������������       �               H�4H�4@������������������������       �      �<       ��/���@�       �                  ;��?�����?       p�[50@������������������������       �               �C=�C=@�       �                 �+�[?"1����?       �`O��"@�       �                 �fQ?;�N9���?       ��{j�@�       �                 pa��?b,���O�?       ���/>@������������������������       �               ��#���?������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?������������������������       �      ��       0#0#@�       �                  �9��?�-l�Fb�?       vrgN�3=@�       �                 ���?�J���?       ��*]Y@������������������������       �               ��#�� @������������������������       �               0#0# @�       �                 p��?t(.�?       Q��9@������������������������       �               %S2%S27@������������������������       �      ȼ       ��/����?�       �                 ���?���߫k�?3       i�ȃ?U@�       �                 ���?$ k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      ��       ��/���@�       �                   ��?�Pq��$�?/       Q� ��T@�       �                 �\�?�9����?!       Km�!�I@�       �                 ��i�?`,�#6?�?
       ���*4@�       �                 ʎ ]?X�ih�<�?       ��
@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                 P���?      �<       ��8��8*@������������������������       �               H�4H�4@������������������������       �               ��+��+$@�       �                 ���?����A��?       ����?@������������������������       �               ��/����?�       �                 �qҍ?RtU���?       �8ܭ�=@�       �                 Ѐ�?|�و��?       cR4��/@�       �                 �� �?���!��?       �@��&@������������������������       �               ��#���?�       �                 ��?Hy��]0�?       ���y"@������������������������       �               ��+��+@������������������������       �      ȼ       ��/����?�       �                 �L��?��^���?       ���w!@�       �                  ��^�?|�G���?       ��%�|@������������������������       �      �<       ��/����?������������������������       �               0#0# @������������������������       �               0����/@������������������������       �        
       �C=�C=,@�       �                 �D�����԰?       �����0<@�       �                 @�P�?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      ��       k�6k�69@�t�bh�hhK ��h��R�(KK�KK��h �B8  U^Cyc@0����/c@� � �d@YUUUU5a@�e�_��W@;�;�F@���>��\@h
��V@��-��-5@w�}w\@鰑U@��8��8*@�k(���U@������S@#0#0&@��,���Q@��h
�G@H�4H�4@�k(���5@�_��e�=@0#0# @������3@��/���.@0#0# @������3@鰑%@        �k(��2@0����/@        �k(��2@��/���@        ��b:��*@��/���@        �k(��"@                ��#��@��/���@                ��/���@        ��#��@                ;��,��@                        ��/����?        ��#���?�cp>@                �cp>@        ��#���?                        0����/@0#0# @        0����/@                        0#0# @��#�� @��|��,@                0����/#@        ��#�� @0����/@        ��#�� @��/����?                ��/����?        ��#�� @                        �cp>@        6��tSH@D�JԮD1@0#0#@6��tSH@��/���.@0#0#@���#8E@���-��@0#0# @���b:@@��/����?        z�5��@��/����?        ;��,��@                ��#���?��/����?        ��#���?                        ��/����?        �#���9@                <��,��$@0����/@0#0# @��#���?0����/@0#0# @        0����/@        ��#���?        0#0# @��#���?                                0#0# @�k(��"@                z�5��@D�JԮD!@0#0# @z�5��@D�JԮD!@        ��#�� @��/����?        ��#�� @                        ��/����?        ��#���?��/���@        ��#���?��/����?                ��/����?        ��#���?                        �cp>@        z�5��@        0#0# @z�5��@                                0#0# @        ��/����?        ��#��0@�]�ڕ�?@��+��+@\Lg1��&@0����/#@        ;��,��$@0����/@        ;��,��@0����/@        ��#��@��/����?                ��/����?        ��#��@                ��#�� @                ��#�� @                ��#���?��/���@                �cp>@        ��#���?��/����?        ��#���?                        ��/����?        ;��,��@                ��#���?0����/@        ��#���?                        0����/@        ;��,��@h
��6@��+��+@z�5��@/����/3@0#0#�?        ���-��*@        z�5��@�cp>@0#0#�?z�5��@��/����?                ��/����?        z�5��@                        ��/���@0#0#�?        ��/���@                        0#0#�?��#�� @�cp>@0#0#@        ��/����?        ��#�� @��/����?0#0#@        ��/����?0#0#@                H�4H�4@        ��/����?0#0#�?                0#0#�?        ��/����?        ��#�� @                ��b:��:@�cp>@0#0# @        ��/����?        ��b:��:@��/���@0#0# @��b:��:@��/���@        �k(��"@��/���@        �k(��"@��/����?        z�5��@��/����?        z�5��@                        ��/����?        z�5��@                        ��/����?        ��,���1@                                0#0# @��#�� @��/���@0#0# @��#�� @��/���@��+��+@��#���?��/���@0#0#�?        ��/���@0#0#�?        ��/���@                        0#0#�?��#���?                ��#���?        0#0#@                0#0# @��#���?        0#0# @                0#0# @��#���?                                H�4H�4@�k(���5@��/���@H�4H�48@<��,��$@��/����?0#0#�?        ��/����?        ;��,��$@        0#0#�?�k(��"@                ��#���?        0#0#�?��#���?                                0#0#�?[Lg1��&@���-��@%S2%S27@�k(��"@�cp>@0#0# @��#�� @�cp>@0#0#�?        �cp>@        ��#�� @        0#0#�?��#�� @                                0#0#�?���>��@        0#0#�?���>��@                                0#0#�?��#�� @��/����?��-��-5@        ��/����?��)��)3@        ��/����?�C=�C=@        ��/����?                        �C=�C=@                H�4H�4(@��#�� @        0#0# @                0#0# @��#�� @                ���>��,@��|��L@�A�A^@z�5��(@鰑E@������J@;��,��$@&jW�v%D@�C=�C=<@��#��@�cp>�9@H�4H�4@��#��@�cp>'@H�4H�4@��#���?        0#0# @��#���?                                0#0# @z�5��@�cp>'@0#0#�?z�5��@�cp>'@        ��#���?�cp>'@        ��#���?��/����?        ��#���?                        ��/����?                /����/#@        ��#�� @                                0#0#�?        ��|��,@        z�5��@��|��,@k�6k�69@;��,��@���-��*@#0#0&@                H�4H�4@;��,��@���-��*@0#0# @;��,��@0����/#@0#0# @        ���-��@0#0# @        �cp>@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @        ��/����?                ��/���@        ;��,��@�cp>@        ;��,��@                        �cp>@                ��/���@H�4H�4@                H�4H�4@        ��/���@        ��#���?��/����?�C=�C=,@                �C=�C=@��#���?��/����?�C=�C=@��#���?��/����?H�4H�4@��#���?        H�4H�4@��#���?                                H�4H�4@        ��/����?                        0#0#@��#�� @��/����?k�6k�69@��#�� @        0#0# @��#�� @                                0#0# @        ��/����?%S2%S27@                %S2%S27@        ��/����?        ��#�� @��/���.@J�dJ��P@��#���?��/���@        ��#���?                        ��/���@        ��#���?�cp>'@K�dJ��P@��#���?鰑%@��+��+D@        ��/����?��)��)3@        ��/����?H�4H�4@        ��/����?                        H�4H�4@                ��8��8*@                H�4H�4@                ��+��+$@��#���?0����/#@��-��-5@        ��/����?        ��#���?��/���@��-��-5@��#���?��/���@�C=�C=@��#���?��/����?��+��+@��#���?                        ��/����?��+��+@                ��+��+@        ��/����?                ���-��@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @        0����/@                        �C=�C=,@        ��/����?�;�;;@        ��/����?0#0# @        ��/����?                        0#0# @                k�6k�69@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ���bhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKυ�h��BH-         �                 p��{?47�LJ�?"      �8��Gs}@       �                 �WR�?p&�C��?�       G"0��w@       p                 ��??<_����?�       	�=o��r@       ?                    �?`��C���?�       ��ډ�j@       $                 )DW?Լ��9��?O       �M���^@       !                 �#h?,=؇��?)       r�go'P@                        �U��������?'       �h�d��N@                        �I?�\�sF��?       U>��1@	                        0��?ދA&w(�?
       �]��0@
                        P���>�����?       ��X�)B @                        @.��>l%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ;��,��@                        �L�^?>ǵ3���?       �q�ͨ�@������������������������       �               ��/���@                       �@B_?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@������������������������       �               ��#���?                          E(�?���+@�?       ���
$F@                         \�&?BF�X��?       -�=k�U0@                         ��G�?���/��?       @z$S��@                         �q�?�����?       ��X�)B@                        �a?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �      м       ��/����?������������������������       �      ȼ       <��,��$@                          U��>      �<       *�����;@������������������������       �               z�5��@������������������������       �               z�5��8@"       #                  �9��?dn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @%       >                 �h�?JO=x��?&       E�_�B�K@&       3                 � l?e������?#       nAw�gJ@'       0                  �q�?t	���?       r�o�`?@(       /                   E(�?rf�T6|�?       x,*��P;@)       .                 .w�S?���/��?       @z$S��'@*       -                 P��r?`n����?       ~��Y-"@+       ,                 �)88?4=�%�?       �(J��@������������������������       �               ��#�� @������������������������       �               �cp>@������������������������       �               ��#��@������������������������       �      Լ       �cp>@������������������������       �      ��	       ��/���.@1       2                 �۶�?f,���O�?       ���/>@������������������������       �               H�4H�4@������������������������       �               ��#���?4       ;                  ��^�?ģ�cE��?       b�co5@5       8                  �9��?�b8�Y�?       HJͰ(@6       7                 `���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?9       :                 ��`?      �<	       <��,��$@������������������������       �               ��#���?������������������������       �               �k(��"@<       =                   ��?Rn����?       ~��Y-"@������������������������       �               �cp>@������������������������       �      ��       z�5��@������������������������       �               z�5��@@       [                 �s��?�b���N�?4       ���JW@A       X                 �;�?���"���?!       �_�q�~O@B       G                 p��?n��H��?       U'y�LH@C       F                 �ĉp?����?       �Ä�>c(@D       E                 �$I�?�)z� ��?       �\�@������������������������       �               �cp>@������������������������       �               ��#��@������������������������       �      ��       ;��,��@H       S                 ��%~?�XӐ���?       \�W=�3B@I       J                hC�Z8?FG�:">�?       �K��G:@������������������������       �               ��#���?K       R                 �Us9?�L����?       [k���>9@L       M                 `��?<f��x��?       Ɋm68@������������������������       �      м
       D�JԮD1@N       Q                  ���?r��H��?       v�I�@O       P                 X��u?����?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?������������������������       �               �cp>@������������������������       �      �<       ��#���?T       U                 пv�?tP�D�?       �A��P?$@������������������������       �               ��#��@V       W                  @V��?���/��?       @z$S��@������������������������       �               z�5��@������������������������       �               �cp>@Y       Z                  �j?      �<       ��|��,@������������������������       �               ��On�(@������������������������       �               ��/����?\       g                 �C�?D�	4�?       ��ߺ4=@]       `                 �Q��?��A=d'�?
       k'��.@^       _                ���ms?      �<       <��,��$@������������������������       �               z�5��@������������������������       �               ��#��@a       f                 ���?:�N9���?       ��{j�@b       e                 `F�?f,���O�?       ���/>@c       d                 е?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �      ȼ       ��/����?h       o                 �ڡ3?�Z�ܙ�?	       c����+@i       j                   .p�?���mf�?       寠�?b#@������������������������       �               ��/���@k       n                  L۰?�� ��?       rp� k@l       m                 ��=�?���mf�?       毠�?b@������������������������       �      �<       ��/���@������������������������       �               0#0#�?������������������������       �               0#0#�?������������������������       �               ��#��@q       �                 p&�?�{%�?7       ���b�V@r       �                  �_�?�*I���?4       ~>�$�U@s       x                  �x��?֙�P�?,       �,�<HR@t       w                 ��I?P���J��?       ��k(/D@u       v                  ;��?$ k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?������������������������       �               ����z�A@y       �                  � �?H^�ZK�?       ���Qa@@z       {                 @F��)�����?       
�p[C1@������������������������       �               z�5��@|       }                 �z�?�����?       W!��&@������������������������       �               �cp>@~       �                 (��?�J���?       ��*]Y @       �                   �0�?�o���?       o�9�F@������������������������       �               ��#���?������������������������       �               0#0#@������������������������       �               z�5��@�       �                   Y��?JW���?
       �$!��.@�       �                 '4�h?@��~d��?	       6E���*@������������������������       �               E�JԮD!@�       �                 h�լ?���mf�?       毠�?b@������������������������       �               0#0#�?������������������������       �      �<       ��/���@������������������������       �               0#0# @�       �                  �0��?�PJo�x�?       T|qt�&@������������������������       �               z�5��@�       �                 ���?:ǵ3���?       �q�ͨ�@������������������������       �               z�5��@�       �                  x\�?      �<       0����/@������������������������       �               ��/����?������������������������       �               ��/���@�       �                 �؉�?E#���?       �B�j@������������������������       �               0#0#@������������������������       �               ��#�� @�       �                 �'f�?U��,��?0       �H�'=�R@�       �                 �vQ?�	J���?(       ��WtuaN@�       �                  �x��?�X�?       n]�
x=@�       �                 �Q�?d%@�"�?       ��[�@�       �                 �r�?$ k�Lj�?       �q��l}@������������������������       �      �<       ��/���@������������������������       �               ��#���?������������������������       �               ��#���?�       �                 0�rM?�}����?       w��H!7@�       �                 0�2�?�IQ���?       ��]4@�       �                    �?��]�uJ�?       ���:O.@�       �                 ��?�k��?       �0QqX@�       �                 ����?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?������������������������       �               0#0#@������������������������       �               0#0# @�       �                  �0��?hutee�?       Q9��@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                 KL�?��q�R�?       C}Ԥ@������������������������       �               ��#���?�       �                 p�'�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 �'Q�?�}h��?       ���r�?@�       �                 ���?��N�O��?       =T�8�2@�       �                 p$�?� �_rK�?       J�@��"@������������������������       �               ��/����?�       �                 ���x?�_�A�?       肵�e`@������������������������       �               ��/����?������������������������       �               ;��,��@�       �                 `�	�?      �<       0����/#@������������������������       �               �cp>@������������������������       �               ���-��@�       �                  ���?P�#O���?       �wtJ*@�       �                 �qp�?�o���?       o�9�F@�       �                 ʊ�X?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               H�4H�4@�       �                 �^��?r�T���?       ��e[�& @������������������������       �               ��#�� @�       �                  ��^�?��q�R�?       B}Ԥ@������������������������       �               ��#�� @�       �                 Pj��?x�G���?       ��%�|@������������������������       �               0#0#�?�       �                  `%+�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                  Ц6�?x��ճC�?       y��l$,@�       �                    �?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               #0#0&@�       �                 `I9�?��4sր�?8       OZ4miW@�       �                 @��?����|e�?       8\@��'@������������������������       �               vb'vb'"@������������������������       �      �<       �cp>@������������������������       �        2       �N��NlT@�t�b��     h�hhK ��h��R�(KK�KK��h �Bh  g:��,&c@�H��tXe@���~�gb@g:��,&c@;�œ[�d@�C=�C=L@k1��tVa@\<�œb@��)��)3@+���>�]@�H��tXU@0#0# @�YLgqT@����z�A@H�4H�4@��b:��J@鰑%@        �#���I@0����/#@        <��,��$@���-��@        �k(��"@���-��@        z�5��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ;��,��@                z�5��@0����/@                ��/���@        z�5��@��/����?                ��/����?        z�5��@                ��#���?                >��,��D@�cp>@        ��b:��*@�cp>@        z�5��@�cp>@        z�5��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                        ��/����?        <��,��$@                *�����;@                z�5��@                z�5��8@                ��#�� @��/����?                ��/����?        ��#�� @                ,�����;@��On�8@H�4H�4@|�5��8@��On�8@H�4H�4@���>��@鰑5@H�4H�4@z�5��@鰑5@        z�5��@�cp>@        z�5��@�cp>@        ��#�� @�cp>@        ��#�� @                        �cp>@        ��#��@                        �cp>@                ��/���.@        ��#���?        H�4H�4@                H�4H�4@��#���?                ��,���1@��/���@        \Lg1��&@��/����?        ��#���?��/����?                ��/����?        ��#���?                <��,��$@                ��#���?                �k(��"@                z�5��@�cp>@                �cp>@        z�5��@                z�5��@                �k(��B@��On�H@��+��+@�k(���5@�)�B�D@        �k(���5@���-��:@        �k(��"@�cp>@        ��#��@�cp>@                �cp>@        ��#��@                ;��,��@                z�5��(@�e�_��7@        ;��,��@鰑5@        ��#���?                ��#��@鰑5@        z�5��@鰑5@                D�JԮD1@        z�5��@��/���@        z�5��@��/����?        z�5��@                        ��/����?                �cp>@        ��#���?                ���>��@�cp>@        ��#��@                z�5��@�cp>@        z�5��@                        �cp>@                ��|��,@                ��On�(@                ��/����?        �P^Cy/@D�JԮD!@��+��+@[Lg1��&@��/����?H�4H�4@<��,��$@                z�5��@                ��#��@                ��#���?��/����?H�4H�4@��#���?        H�4H�4@��#���?        0#0#�?                0#0#�?��#���?                                0#0# @        ��/����?        ��#��@��/���@0#0# @        ��/���@0#0# @        ��/���@                ��/���@0#0# @        ��/���@0#0#�?        ��/���@                        0#0#�?                0#0#�?��#��@                ������3@�_��e�M@#0#0&@��,���1@�_��e�M@�C=�C=@ZLg1��&@\�v%jWK@�C=�C=@��#���?������C@        ��#���?��/���@                ��/���@        ��#���?                        ����z�A@        <��,��$@��/���.@�C=�C=@<��,��$@�cp>@0#0#@z�5��@                ��#��@�cp>@0#0#@        �cp>@        ��#��@        0#0#@��#���?        0#0#@��#���?                                0#0#@z�5��@                        ��On�(@H�4H�4@        ��On�(@0#0#�?        E�JԮD!@                ��/���@0#0#�?                0#0#�?        ��/���@                        0#0# @z�5��@0����/@        z�5��@                z�5��@0����/@        z�5��@                        0����/@                ��/����?                ��/���@        ��#�� @        0#0#@                0#0#@��#�� @                ���>��,@�cp>7@�z��z�B@���>��,@h
��6@H�4H�48@��#��@���-��@vb'vb'2@��#�� @��/���@        ��#���?��/���@                ��/���@        ��#���?                ��#���?                ��#�� @�cp>@vb'vb'2@��#���?��/����?S2%S2%1@��#���?        �C=�C=,@��#���?        H�4H�4@��#���?        0#0# @                0#0# @��#���?                                0#0#@                0#0# @        ��/����?H�4H�4@        ��/����?                        H�4H�4@��#���?��/����?0#0#�?��#���?                        ��/����?0#0#�?        ��/����?                        0#0#�?;��,��$@��/���.@H�4H�4@;��,��@���-��*@        ;��,��@��/���@                ��/����?        ;��,��@��/����?                ��/����?        ;��,��@                        0����/#@                �cp>@                ���-��@        ;��,��@��/����?H�4H�4@��#���?        0#0#@��#���?        0#0#�?��#���?                                0#0#�?                H�4H�4@��#��@��/����?0#0# @��#�� @                ��#�� @��/����?0#0# @��#�� @                        ��/����?0#0# @                0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                ��/����?��8��8*@        ��/����?0#0# @        ��/����?                        0#0# @                #0#0&@        �cp>@;�;�V@        �cp>@vb'vb'"@                vb'vb'"@        �cp>@                        �N��NlT@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ+�MhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK煔h��B�2         x                    �?D���Q�?!      ���*5�}@       ;                 ����?������?�       &P@�}m@       (                 �)�4?tt2pY�?@       g��L/�Z@       #                 �@�?2�@��?,       �8����R@                        `��u?Ga�]��?(       x��G�P@                        �+"�?<Bms�?        ��֖��K@                        x��?X�:V��?       �K��GJ@                        �L'?M�����?       q����.@	                        �^&?��t� �?	       ����x&@
                        P���>      �<       z�5��@������������������������       �               ��#���?������������������������       �               ;��,��@                         Ц6�?ܗZ�	7�?       j~���@                         �G?�?f%@�"�?       ��[�@������������������������       �               ��/����?                        &H�9?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �      м       ��#��@                        P�y?��p?��?       P�^��B@                         �]m?d�s�	�?       f���*@������������������������       �               ��/����?������������������������       �               z�5��(@������������������������       �      �<       �,����7@                        P��?dn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @                        Ĕ~?�����?       �Ä�>c(@������������������������       �               ��/����?       "                 ��s?��t� �?       ����x&@        !                ����?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#�� @$       '                 GW�d?�LU���?       i�ҹ^�@%       &                  ���?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �               ��/���@)       4                  s��?9B���M�?       ߒ��F�>@*       1                 ��M�?f�4��d�?       ,�V��v3@+       0                 P>-l?r@ȱ��?       ���~1@,       -                 ��?�h��%�?
       �1�
�u0@������������������������       �               0����/#@.       /                 �\�?��|��?       ���ĺw@������������������������       �               0����/@������������������������       �               ��#�� @������������������������       �      �<       ��#���?2       3                 ���?��G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?5       6                  �`<?�cj����?       f�e�JO&@������������������������       �               ��/����?7       :                 @��?X����1�?       �����x"@8       9                `?�j�?b,���O�?       ���/>@������������������������       �               ��#���?������������������������       �               H�4H�4@������������������������       �               ;��,��@<       u                 ��g?������?V       t���v9`@=       r                 �Fܴ?�w��#�?:       k}�g�U@>       i                 0�?v֥�3��?7       �y��]�T@?       \                  �/�?D���Rg�?.       焙��P@@       S                 `���?�%#���?       ���JE@A       R                  @���?�=vo�`�?       �M��Jg?@B       C                 �i�N?����?       ��.�SU=@������������������������       �               z�5��@D       I                 �\ͥ?*��_ H�?       �q^a::@E       H                 p
I�?���`�?       ��
�Me@F       G                 @+{�?r@ȱ��?       om���S@������������������������       �               0����/@������������������������       �               ��#���?������������������������       �               0#0# @J       Q                   ��?��%�U��?       o/o�a2@K       L                 �lY�?2 k�Lj�?       �q��l}#@������������������������       �               �cp>@M       P                 �Ӝ�?���/��?       V��7�@N       O                 p��!?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      �<       ��/����?������������������������       �               E�JԮD!@������������������������       �      �<       ��#�� @T       W                   E(�?�"�F��?
       >�h�\&@U       V                ��F�u?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?X       [                 ����?x�t1u�?       "�te!� @Y       Z                 ��aӾ�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �      ��       z�5��@]       d                 �m�?J=W���?       �CJ��^9@^       c                �s�t?8�s�	�?	       f���*@_       b                 x�g�?�����?       �O��@`       a                 p�M�?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               z�5��@������������������������       �      �<       ���>��@e       h                 H�	�?�\U�?       �{����'@f       g                  �{��?��[����?       Hl�_A@������������������������       �               0����/@������������������������       �               0#0# @������������������������       �               ;��,��@j       o                 @Ws�?d9����?	       }��.�,@k       l                 ���@?�+�z���?       KGh��
)@������������������������       �      ��       E�JԮD!@m       n                 @�C�?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@p       q                  0Y��?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?s       t                  p��?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@v       w                 �@A�?      �<       �
��
�E@������������������������       �               0#0# @������������������������       �               �ڬ�ڬD@y       �                  �g<�?&������?�       se�ܔm@z       �                 `*X�?Jry���?*       sm�S@{       �                  �?��{@��?       ��I�@B@|       �                 p�%c?�Ug���?       ����0@}       �                 P��?^%@�"�?       ��[�'@~                        p�R?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @�       �                 ���B?fQ��?       �s�=�!@������������������������       �               ��#���?�       �                  h��?`�r{��?       e�6� @�       �                 ���\?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �               0����/@������������������������       �      �<       ;��,��@�       �                 �=�?@#����?       w�߄�3@������������������������       �               ;��,��$@�       �                 �M��?D���'0�?       �C�� T"@������������������������       �               ��#��@�       �                 ��?��Z�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@�       �                 ą�s?�̥Q)�?       �F�C@�       �                 ˢ?������?       jƹ�J�;@�       �                �s�[w?��oR��?       m�Q6�(@�       �                 ���?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      �<       ;��,��$@�       �                  �?pLU���?
       h�ҹ^�.@������������������������       �        	       ���-��*@������������������������       �               0#0# @������������������������       �      ȼ       H�4H�4(@�       �                 Фͽ?��^r��?a       ��=�d@�       �                 x�	�?-��?'       �0�?P@�       �                  `K�?���H��?"       ���|��K@�       �                 ��x�?�p�Nt�?       ����C@�       �                 �j��?���d���?       zu��A@�       �                 ���?,��hz��?       �
�j9@�       �                 ��s?��oB��?       ���m2@�       �                 �/?�(���?       y��uk1@�       �                 �[l?, k�Lj�?       �q��l}#@������������������������       �               ��/���@�       �                 @�>b%@�"�?       ��[�@������������������������       �      �<       ��/���@������������������������       �               ��#�� @������������������������       �      ��       ��/���@������������������������       �               0#0#�?�       �                 0��?���1p8�?       |곯�@������������������������       �               0#0#@�       �                   ��?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 @�V?      �<       鰑%@������������������������       �               ��/����?������������������������       �               D�JԮD!@�       �                   �0�?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?�       �                 �j��?jn����?       Ҁh��K.@������������������������       �               z�5��@�       �                 ����?��<��?
       s=�x�(@�       �                  ��?@���'0�?       �C�� T"@�       �                 d���?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                  �!�?\����?       P	K��@������������������������       �               ��/����?������������������������       �               z�5��@������������������������       �      Լ       �cp>@�       �                  �Ԧ�?jutee�?       Q9��#@������������������������       �               H�4H�4@�       �                 @��?�w��d��?       �0���s@������������������������       �      �<       H�4H�4@������������������������       �               ��/���@�       �                 0�=�?H�|g�?:       œ���W@�       �                 ���?Rہ(J�?-       �Z��CQ@�       �                 ��j�?���j��?%       �X���L@�       �                 Ќ�j? �
Fq�?       /��C@�       �                 ���?@˒�0�?       �A��Z!5@�       �                  �g�?����|e�?       �z �B�@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?������������������������       �      ��	       S2%S2%1@�       �                 p.�?:�4��?       p��P9�0@�       �                 � ��?�n���k�?	       3��&�*@������������������������       �               vb'vb'"@�       �                 �I�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �      ȼ       ��/���@�       �                 p���?\�}R4�?       �[RZ��3@�       �                 CJ�?J5�,�r�?	       7�r|k\,@�       �                 7�?�4^��?       s_w$/"@�       �                 8��?���/��?       V��7�@������������������������       �               ��/����?�       �                  L�?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               ��+��+@�       �                 p��?L� P?)�?       ����x�@������������������������       �               0#0#�?������������������������       �               ��#��@�       �                 �!�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/���@�       �                 �+�[?      �<       #0#0&@������������������������       �               ��+��+@������������������������       �               H�4H�4@������������������������       �      ��       ��8��8:@�t�bh�hhK ��h��R�(KK�KK��h �B�  	��GPd@��e�_�b@��+��+d@�#���Y@;l��F:R@����M@��,���Q@��/���>@��+��+@��>���N@���-��*@0#0#�?��>���N@���-��@        �#���I@��/���@        |�5��H@�cp>@        ��b:��*@��/����?        �k(��"@��/����?        z�5��@                ��#���?                ;��,��@                z�5��@��/����?        ��#���?��/����?                ��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#�� @                ��#��@                �YLg1B@��/����?        {�5��(@��/����?                ��/����?        z�5��(@                �,����7@                ��#�� @��/����?                ��/����?        ��#�� @                �k(��"@�cp>@                ��/����?        �k(��"@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                        ���-��@0#0#�?        �cp>@0#0#�?                0#0#�?        �cp>@                ��/���@        �k(��"@D�JԮD1@0#0#@z�5��@��/���.@0#0#�?z�5��@��|��,@        ��#�� @��|��,@                0����/#@        ��#�� @0����/@                0����/@        ��#�� @                ��#���?                        ��/����?0#0#�?        ��/����?                        0#0#�?z�5��@��/����?H�4H�4@        ��/����?        z�5��@        H�4H�4@��#���?        H�4H�4@��#���?                                H�4H�4@;��,��@                ��#��@@鰑E@�;�;K@��#��@@鰑E@#0#0&@��#��@@�)�B�D@0#0# @��#��@@��|��<@H�4H�4@�P^Cy/@�cp>7@0#0#@��#�� @鰑5@0#0# @z�5��@鰑5@0#0# @z�5��@                z�5��@鰑5@0#0# @��#���?0����/@0#0# @��#���?0����/@                0����/@        ��#���?                                0#0# @��#�� @Nn��O0@        ��#�� @��/���@                �cp>@        ��#�� @��/����?        ��#�� @��/����?        ��#�� @                        ��/����?                ��/����?                E�JԮD!@        ��#�� @                ���>��@��/����?0#0# @        ��/����?0#0#�?                0#0#�?        ��/����?        ���>��@        0#0#�?��#���?        0#0#�?                0#0#�?��#���?                z�5��@                ��,���1@�cp>@0#0# @z�5��(@��/����?        ;��,��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        z�5��@                ���>��@                ;��,��@0����/@0#0# @        0����/@0#0# @        0����/@                        0#0# @;��,��@                        ��On�(@0#0# @        �cp>'@0#0#�?        E�JԮD!@                �cp>@0#0#�?                0#0#�?        �cp>@                ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?H�4H�4@        ��/����?                        H�4H�4@                �
��
�E@                0#0# @                �ڬ�ڬD@    �M@v�'�x�R@w?�s?wY@�k(��B@�e�_��7@�A�A.@��b:��:@/����/#@        �k(��"@��/���@        ��#��@��/���@        ��#�� @��/����?                ��/����?        ��#�� @                ��#�� @���-��@        ��#���?                ��#���?���-��@        ��#���?��/����?                ��/����?        ��#���?                        0����/@        ;��,��@                ��,���1@��/����?        ;��,��$@                ���>��@��/����?        ��#��@                z�5��@��/����?                ��/����?        z�5��@                ;��,��$@��|��,@�A�A.@;��,��$@��|��,@H�4H�4@;��,��$@��/����?0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?;��,��$@                        ���-��*@0#0# @        ���-��*@                        0#0# @                H�4H�4(@�k(���5@�cp>�I@�
��
�U@�P^Cy/@0����/C@#0#0&@�P^Cy/@F�JԮDA@��+��+@;��,��@�_��e�=@��+��+@z�5��@�a#6�;@��+��+@z�5��@D�JԮD1@��+��+@��#�� @��/���.@0#0#�?��#�� @��/���.@        ��#�� @��/���@                ��/���@        ��#�� @��/���@                ��/���@        ��#�� @                        ��/���@                        0#0#�?��#���?��/����?0#0#@                0#0#@��#���?��/����?        ��#���?                        ��/����?                鰑%@                ��/����?                D�JԮD!@        ��#�� @��/����?        ��#�� @                        ��/����?        <��,��$@0����/@        z�5��@                ���>��@0����/@        ���>��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        z�5��@��/����?                ��/����?        z�5��@                        �cp>@                ��/���@H�4H�4@                H�4H�4@        ��/���@H�4H�4@                H�4H�4@        ��/���@        z�5��@���-��*@�i��R@z�5��@���-��*@]��Y��H@z�5��@���-��*@��)��)C@        �cp>@0#0#@@        ��/����?��+��+4@        ��/����?H�4H�4@                H�4H�4@        ��/����?                        S2%S2%1@        0����/@H�4H�4(@        ��/����?H�4H�4(@                vb'vb'"@        ��/����?H�4H�4@        ��/����?                        H�4H�4@        ��/���@        z�5��@��/���@H�4H�4@z�5��@��/����?H�4H�4@��#�� @��/����?��+��+@��#�� @��/����?                ��/����?        ��#�� @��/����?        ��#�� @                        ��/����?                        ��+��+@��#��@        0#0#�?                0#0#�?��#��@                        �cp>@                ��/����?                ��/���@                        #0#0&@                ��+��+@                H�4H�4@                ��8��8:@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJY]hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKх�h��B�-         T                 �'��?��տO�?&      H�;�}@       5                  ����?���Rx��?|       ��Q�h@       (                 �l�A?�t�A��?H       W��*�\@       	                 �@?(�0�7�?2       � %��S@                        ��V?��t� �?       ����x6@                        ��IL?� �_rK�?       J�@��"@������������������������       �               ;��,��@������������������������       �      ��       ��/���@������������������������       �        	       ��b:��*@
                        ���D?@H�o�?#       ���D�K@������������������������       �               0����/@                        �
ǂ?#].��?!       {˸ II@                        @*��? Z��K�?       ��K�M�:@                        �K?�_�A�?	       肵�e`,@������������������������       �               ��#��@                        @�?��Z�	7�?       i~���$@                        hf�?����?       ��X�)B @������������������������       �               ��/����?                         @mj�?l����?       P	K��@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?                         @(B�?,��c`�?       %��t5)@                           �?      �<       0����/#@������������������������       �               ��/���@������������������������       �               �cp>@                       ��}Ez?^%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?       '                  s��?T�1�7�?       l&sDB8@                         @���?�������?       ���|a5@������������������������       �               |�5��(@!       &                 8��?`���?       ��Me�!@"       %                  �9��?j��H��?       v�I�@#       $                 (b�q?$ k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      ��       ��/���@������������������������       �               ��#�� @������������������������       �               0#0# @������������������������       �      �<       �cp>@)       ,                  �0��?D��M�?       6B��	�B@*       +                 @F��d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@-       2                 е�?8*9��?       9��g��?@.       /                  �"�?0\qi�H�?       ��%@f�<@������������������������       �        
       ��/���.@0       1                 �S�?D��~d��?       8E���*@������������������������       �               ��On�(@������������������������       �               0#0#�?3       4                    �?H����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?6       Q                  k��?f���W�?4       	����T@7       N                 �f�V?җ��?0       +�E�i[S@8       K                 �y����my����?,       M���H$Q@9       H                 �� �?��C����?       �o>��,7@:       E                   p��?&��˕j�?       �q�ހA5@;       B                    �?֥��Y��?       �u%!!k1@<       ?                 �Z�?�.��8��?       �,_�.@=       >                 ��x�?����X��?       &��֞&@������������������������       �               ;��,��$@������������������������       �      ȼ       ��/����?@       A                 ��a�?�zœ���?       IG���t@������������������������       �               z�5��@������������������������       �               0#0#�?C       D                 @��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?F       G                 .25Q?      �<       ��/���@������������������������       �               �cp>@������������������������       �               ��/����?I       J                    �?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?L       M                 `�?�(1k��?       �ꁞ9�F@������������������������       �               �k(���E@������������������������       �      �<       ��/����?O       P                  䈂?z%@�"�?       �6�E�!@������������������������       �               �cp>@������������������������       �      ȼ       z�5��@R       S                 �� �?�@����?       ���a�@������������������������       �               ��/����?������������������������       �               0#0#@U       �                 ���?�=�4�8�?�       ��Ȓ�'q@V       �                 ��@s?՜��-��?�       {k�[(j@W       �                 ��K?u�x!m��?Y       Kŏa@X       {                 ���s?�<��?�?A       3���c�Y@Y       x                  ��?f�/W�D�?$       ,�.�@K@Z       u                 ��x�?憛���?!       �őSA�H@[       \                  L��?R�H�q�?       pM��$F@������������������������       �               H�4H�4@]       h                 @��?�-*����?       :�ǀ�D@^       g                 wȧ?BW���?
       �$!��.@_       d                 �J�?x9����?	       |��.�,@`       a                 ��gn?�@G���?       hu��@������������������������       �               �cp>@b       c                 `U�?h�4���?       �tCP��@������������������������       �               0#0# @������������������������       �               �cp>@e       f                 �k��?      �<       ���-��@������������������������       �               ��/����?������������������������       �               0����/@������������������������       �               0#0#�?i       n                  ��?ࢡF$Y�?       �����9@j       m                 Е��?�`@s'��?
       Di_y,*+@k       l                 �U��>`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               鰑%@o       t                    �?b,���O�?	       ԥ��G](@p       s                 �p��?�ctn�0�?       �$�k�K @q       r                  ;��?�zœ���?       IG���t@������������������������       �               0#0#�?������������������������       �               z�5��@������������������������       �      ��       0#0#@������������������������       �               0#0#@v       w                 ���?      �<       ��+��+@������������������������       �               0#0#�?������������������������       �               0#0#@y       z                   E(�?      �<       ;��,��@������������������������       �               ��#�� @������������������������       �               z�5��@|       �                 �3��?O��Z*�?       :��H@}       �                 F'�?���AK�?       _I��#�B@~       �                    �?��]��?       �nF�f1>@       �                      ��t� �?       ����x&@�       �                 �?      �<       �k(��"@������������������������       �               z�5��@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?�       �                 ����?������?       Ӌ]!_�2@������������������������       �               ��#��@�       �                  �6�?jy�|�?	       (�0�-@�       �                 ��ߢ?�djH�E�?       ^�\m�n@������������������������       �               ��#��@�       �                 0�k�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 ����?)���?       y��uk!@������������������������       �               ���-��@�       �                 �0��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ���>��@�       �                 xb'�?Hj��w�?       l8�(@�       �                  @V��?D��NV=�?       �t�ܲ@������������������������       �               ��#���?�       �                 �Ψ?�� ��?       rp� k@������������������������       �               ��/����?�       �                 0!i�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0# @�       �                 ��?�,�����?       �#$w@@�       �                 ��{�?�1A�]�?       ag	��?@�       �                 h�R?�~�&��?       ?�]��@�       �                 ��j?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �               0#0#@�       �                  �u��? NU�w�?       ���6:&7@�       �                 p���?��/Ѷ?       ���
$6@�       �                  ���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 �}*�?      �<       %jW�v%4@������������������������       �               ��/����?������������������������       �               /����/3@������������������������       �               0#0#�?������������������������       �      �<       ��#���?�       �                 ����?��B��?'       �_�
�KR@�       �                  �E�?Dr����?&       ^����Q@�       �                 �+�[?To��?�?       �>���~C@������������������������       �               ��/����?�       �                 �qҍ?�i\%���?       �����B@�       �                    �?�AP�9��?       h��6��+@������������������������       �               H�4H�4@�       �                 ��?x�G���?       ��%�|@�       �                 �i��?�@����?       ���a�@�       �                  w}?z��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               0#0# @������������������������       �               �cp>@�       �                 �֠�?@4�+W�?       ����%7@�       �                 ��]�?�v�;B��?       ՟���	 @������������������������       �               �C=�C=@������������������������       �      ȼ       ��/����?������������������������       �      �<       �A�A.@������������������������       �               0#0#@@������������������������       �      �<       ��/����?�       �                 `��?p��C 8�?*       E�K�6OP@�       �                 p&�?b� �?       �l��0@�       �                 �x��?���MF�?	       �`�I-*@�       �                 x嶹? v=���?       � ��R(@������������������������       �               ��/����?������������������������       �               #0#0&@������������������������       �      ܼ       ��#���?������������������������       �      ȼ       ��/���@�       �                 �;�?x��fņ�?       ҋ�'H@�       �                  (��?�^�F�M�?       ��ޚ�6@������������������������       �               ��/����?�       �                 P�,�?@˒�0�?       �A��Z!5@������������������������       �      ��       0#0#0@�       �                �톟�?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?������������������������       �               ��8��8:@�t�bh�hhK ��h��R�(KK�KK��h �B�  g:��,&c@q�'�x�b@�fm�f�d@Rg1��4\@s�'�x�R@vb'vb'"@�#���I@�_��e�M@0#0#@]Lg1��F@��/���>@0#0# @�k(��2@��/���@        ;��,��@��/���@        ;��,��@                        ��/���@        ��b:��*@                ��b:��:@���-��:@0#0# @        0����/@        ��b:��:@h
��6@0#0# @ZLg1��&@��/���.@        ;��,��$@��/���@        ��#��@                z�5��@��/���@        z�5��@��/����?                ��/����?        z�5��@��/����?        z�5��@                        ��/����?                ��/����?        ��#���?�cp>'@                0����/#@                ��/���@                �cp>@        ��#���?��/����?                ��/����?        ��#���?                �P^Cy/@���-��@0#0# @�P^Cy/@��/���@0#0# @|�5��(@                z�5��@��/���@0#0# @z�5��@��/���@        ��#���?��/���@        ��#���?                        ��/���@        ��#�� @                                0#0# @        �cp>@        z�5��@��|��<@0#0# @��#��@��/����?                ��/����?        ��#��@                ��#�� @�a#6�;@0#0# @        �a#6�;@0#0#�?        ��/���.@                ��On�(@0#0#�?        ��On�(@                        0#0#�?��#�� @        0#0#�?��#�� @                                0#0#�?��>���N@On��O0@��+��+@��>���N@��/���.@0#0#�?���>��L@0����/#@0#0#�?���>��,@��/���@0#0#�?���>��,@�cp>@0#0#�?���>��,@��/����?0#0#�?��b:��*@��/����?0#0#�?;��,��$@��/����?        ;��,��$@                        ��/����?        z�5��@        0#0#�?z�5��@                                0#0#�?��#���?��/����?        ��#���?                        ��/����?                ��/���@                �cp>@                ��/����?                ��/����?                ��/����?                ��/����?        �k(���E@��/����?        �k(���E@                        ��/����?        z�5��@�cp>@                �cp>@        z�5��@                        ��/����?0#0#@        ��/����?                        0#0#@��k(/D@r�'�x�R@��
���c@������C@F�JԮDQ@o�6k�6Y@������C@=��18N@vb'vb'B@�k(��B@;l��F:B@�A�A>@<��,��$@�e�_��7@��+��+4@;��,��@�e�_��7@��+��+4@;��,��@�e�_��7@�A�A.@                H�4H�4@;��,��@�e�_��7@H�4H�4(@        ��On�(@H�4H�4@        ��On�(@0#0# @        �cp>@0#0# @        �cp>@                �cp>@0#0# @                0#0# @        �cp>@                ���-��@                ��/����?                0����/@                        0#0#�?;��,��@�cp>'@vb'vb'"@��#�� @�cp>'@        ��#�� @��/����?        ��#�� @                        ��/����?                鰑%@        z�5��@        vb'vb'"@z�5��@        ��+��+@z�5��@        0#0#�?                0#0#�?z�5��@                                0#0#@                0#0#@                ��+��+@                0#0#�?                0#0#@;��,��@                ��#�� @                z�5��@                ��b:��:@��On�(@��+��+$@
�#���9@鰑%@0#0#�?�k(��2@鰑%@0#0#�?�k(��"@��/����?        �k(��"@                z�5��@                z�5��@                        ��/����?        �k(��"@E�JԮD!@0#0#�?��#��@                ;��,��@E�JԮD!@0#0#�?��#��@��/����?0#0#�?��#��@                        ��/����?0#0#�?        ��/����?                        0#0#�?��#���?��/���@                ���-��@        ��#���?��/����?        ��#���?                        ��/����?        ���>��@                ��#���?��/����?vb'vb'"@��#���?��/����?0#0#�?��#���?                        ��/����?0#0#�?        ��/����?                ��/����?0#0#�?                0#0#�?        ��/����?                        0#0# @��#�� @�e�_��7@H�4H�4@��#���?�e�_��7@H�4H�4@        �cp>@��+��+@        �cp>@0#0#�?        �cp>@                        0#0#�?                0#0#@��#���?鰑5@0#0#�?��#���?鰑5@        ��#���?��/����?                ��/����?        ��#���?                        %jW�v%4@                ��/����?                /����/3@                        0#0#�?��#���?                        E�JԮD!@1#0#P@        ���-��@0#0#P@        ���-��@0#0#@@        ��/����?                0����/@0#0#@@        ��/���@��+��+$@                H�4H�4@        ��/���@0#0#@        ��/����?0#0#@        ��/����?0#0# @                0#0# @        ��/����?                        0#0# @        �cp>@                ��/����?#0#06@        ��/����?�C=�C=@                �C=�C=@        ��/����?                        �A�A.@                0#0#@@        ��/����?        ��#���?���-��@�[��[�L@��#���?0����/@#0#0&@��#���?��/����?#0#0&@        ��/����?#0#0&@        ��/����?                        #0#0&@��#���?                        ��/���@                ��/����?$S2%S2G@        ��/����?��+��+4@        ��/����?                ��/����?��+��+4@                0#0#0@        ��/����?0#0#@                0#0#@        ��/����?                        ��8��8:@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ4
hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKх�h��B�-         �                 ��{�?[\X?�?(      ��<�}@       �                  �E�?���1�?       ��AĹ�|@       �                 �/��?b����?�       �µE�t@       1                 0-?����l�?�       7�鍅�t@                        `�c?�M:���?8       P����Y@                        �.��?bdؗ��?       4d��8@                        pG�?���.�2�?       ��k	j3@       	                 �-�?f%@�"�?       �6�E�!@������������������������       �               �cp>@
                        `���>      �<       z�5��@������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �      �<       鰑%@                        Z�K?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?       *                  vU{?d�SbA��?(       >�Ҿ�S@                        @��>�x�<�?"       Y&b��qQ@                        ���>���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?       !                 ����?�+op�?        ���ǢrP@                        p�;O?�(1k��?       �ꁞ9�F@                         �P��?�V_�"�?       �����E@������������������������       �        	       �k(���5@                         �Q�?X ����?
       1
C>�5@                           �?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               �k(��2@                         X��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?"       #                 P�?�d�$���?       �T�f4@������������������������       �               ��/����?$       )                 Po?h�j���?
       ���z2@%       &                    �?h�:V��?	       �GP�1@������������������������       �               ZLg1��&@'       (                 �H�=?�����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?������������������������       �      �<       ��/����?+       ,                 ��p?� �_rK�?       J�@��"@������������������������       �               z�5��@-       0                 lj^�?d%@�"�?       ��[�@.       /                ���w?$ k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?������������������������       �               ��#���?2       �                 p��g?F����?�       K�9al@3       f                 ��*?�W#�Z4�?t       ��=g@4       ]                 ��<�?���s��?H       �
!��*]@5       R                 @��?"ϮE�?;       l�
��X@6       7                 �~�X?��#�Jr�?/       +7�'�T@������������������������       �               0����/@8       K                 0S�r?޻��ʫ�?,       xXm")�S@9       J                 ���?4�����?       �W
�ŚA@:       I                 �U��>�uNɗ}�?       S��}@@;       F                  `�J�?���5H�?       ����c9?@<       E                 ��?�?�h�?�C�?       ��=��}6@=       B                 �zz?VB���?       ��>#$$@>       ?                  ��g�?�_�A�?       炵�e`@������������������������       �               ��/����?@       A                 �㐢?�����?       �O��@������������������������       �               ��/����?������������������������       �      �<       ;��,��@C       D                 P��?x��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      �<       z�5��(@G       H                 X���?��^���?       ���w!@������������������������       �               ���-��@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �      �       H�4H�4@L       Q                 `�? �=�Sο?       fY�R��E@M       P                 ��U�?����N-�?       �#[�$E@N       O                 � b?�(߫$��?       0H����*@������������������������       �               ��/����?������������������������       �               [Lg1��&@������������������������       �      �<       ���>��<@������������������������       �      �<       ��/����?S       T                 `��z?p!A_!�?       E����0@������������������������       �               0#0# @U       X                  �Ѱ?��Ik���?       ��c��.-@V       W                  ��d�?�>s{Ab�?       aI��n'@������������������������       �               鰑%@������������������������       �               0#0#�?Y       Z                 ��y�?hn����?       � ��w<@������������������������       �               ��#���?[       \                 `}��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?^       _                    �?P�an41�?       �	Yt�0@������������������������       �               0����/@`       a                 ����?���S&�?	       �3�(@������������������������       �               ��#�� @b       e                 0Y�?&^�yU�?       ��7�1�#@c       d                 �Q�?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �      �<       H�4H�4@g       r                  @mj�?$2$ĝ��?,       �����P@h       i                 Y�b?���:1=�?       ���QE@������������������������       �               ��#�� @j       q                 0*tC?֥�Y��?       %Ճ�HD@k       l                 5��?B��X�&�?       �6��	�@������������������������       �               �cp>@m       n                 ��}�?�nɵ��?       Cad�J@������������������������       �               z�5��@o       p                �6�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               On��O@@s       �                 p��?bYӱA��?       �Nf��8@t       }                  ����?��_�u��?       ��X̰3@u       v                  �~��?H��aB��?       ����"@������������������������       �               0#0#�?w       |                 �38�?@9�)\e�?       _���b @x       {                 ��?�_�A�?       肵�e`@y       z                 P��s?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#��@������������������������       �      м       ��/����?~                        @��?�^�#΀�?       O�{��A%@������������������������       �               D�JԮD!@�       �                   ���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                  ���?�o���?       o�9�F@������������������������       �               0#0#@������������������������       �               ��#���?�       �                  ��^�?�����?       <F"�|E@�       �                 `��?d��Ɵ��?       �(�NA@������������������������       �               ��/����?�       �                 ���?�N�u�?       i���@@�       �                 '4�h?����԰?       �����0<@������������������������       �               ��/����?������������������������       �               �;�;;@�       �                 ��3�?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?�       �                 H��?�����?       �v�qp�!@������������������������       �               0#0#@������������������������       �               0����/@�       �                  p���?      �<       0����/@������������������������       �               ��/����?������������������������       �               �cp>@�       �                   Y��?����?S       ��0��a_@�       �                 p��?��
%��?-       Ӏ���Q@�       �                 v �?:����?       �p�B@�       �                 �ڡC?�:zk���?       �*�]7 ?@�       �                 �@�?>9�)\e�?       ��)8@�       �                    �?�����?       8�nN�R4@�       �                 ���?H�s�	�?	       f���*@������������������������       �               ���>��@�       �                 ��x�?�����?       �O��@������������������������       �               ��/����?������������������������       �      �<       ;��,��@�       �                 @�>t��H��?       v�I�@�       �                  �N�?$ k�Lj�?       �q��l}@������������������������       �               ��/����?�       �                 `��?`%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �      м       ��/���@�       �                 �j'�?��n��?       �-H�\@�       �                 ȍܸ?�֪u�_�?       ��?�8@�       �                  �G?�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               ��+��+@�       �                  �Mm�?�Y�R���?       x��\�A@�       �                    �?w�;B��?       ՟���	@@�       �                 ȯ�?����|e�?
       �z �B�/@������������������������       �               ��/����?�       �                 ��?X�ih�<�?	       ��
,@������������������������       �               ��+��+$@�       �                 lP�w?x�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �        	       0#0#0@�       �                  Q��?x����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @�       �                 |�eO?VN�~��?&       Fi_y,*K@������������������������       �               z�5��@�       �                 ��N�?�\�B7��?"       �Ǣ�9H@�       �                 (�r?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0# @�       �                  �!�?@�z�?       ��B,D@�       �                 ���?     ��?       "F�b@������������������������       �               ��#�� @������������������������       �               H�4H�4@�       �                 ����?��	6?�?       ���J��A@�       �                 pMC�?�^�F�M�?       ��ޚ�&@������������������������       �               ��+��+$@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       H�4H�48@�       �                  ���?�/y߃�?       Ɓ\��((@�       �                 �ɚ�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       ��+��+$@�t�bh�hhK ��h��R�(KK�KK��h �B�       f@P��+c@p�fm��a@�#����e@s�'�x�b@C�A�`@�k(��b@_�_���_@�s?�s?M@�k(��b@��/���^@�s?�s?M@�k(��R@��|��<@        ���>��@D�JԮD1@        z�5��@On��O0@        z�5��@�cp>@                �cp>@        z�5��@                ��#���?                ��#�� @                        鰑%@        ��#��@��/����?        ��#��@                        ��/����?        "�}��P@�cp>'@        �P^CyO@��/���@        ��#�� @��/����?        ��#�� @                        ��/����?        Jp�}N@�cp>@        �k(���E@��/����?        ���#8E@��/����?        �k(���5@                ;��,��4@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        �k(��2@                ��#���?��/����?                ��/����?        ��#���?                ��#��0@��/���@                ��/����?        ��#��0@��/����?        ��#��0@��/����?        ZLg1��&@                ;��,��@��/����?        ;��,��@                        ��/����?                ��/����?        ;��,��@��/���@        z�5��@                ��#�� @��/���@        ��#���?��/���@                ��/���@        ��#���?                ��#���?                �k(��R@~�h
�W@�s?�s?M@�k(��R@��]�ڕU@%S2%S27@�P^CyO@�+Q��B@S2%S2%1@Lp�}N@�_��e�=@��+��+$@���>��L@:l��F:2@�C=�C=@        0����/@        ���>��L@���-��*@�C=�C=@��,���1@鰑%@�C=�C=@��,���1@鰑%@0#0#@��,���1@0����/#@0#0#@��,���1@�cp>@0#0# @;��,��@�cp>@0#0# @;��,��@��/����?                ��/����?        ;��,��@��/����?                ��/����?        ;��,��@                        ��/����?0#0# @        ��/����?                        0#0# @z�5��(@                        ���-��@0#0# @        ���-��@                        0#0# @        ��/����?                        H�4H�4@��k(/D@�cp>@        ��k(/D@��/����?        ZLg1��&@��/����?                ��/����?        [Lg1��&@                ���>��<@                        ��/����?        ��#�� @�cp>'@H�4H�4@                0#0# @��#�� @�cp>'@0#0#�?        鰑%@0#0#�?        鰑%@                        0#0#�?��#�� @��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                ��#�� @��/���@�C=�C=@        0����/@        ��#�� @�cp>@�C=�C=@��#�� @                        �cp>@�C=�C=@        �cp>@0#0#�?                0#0#�?        �cp>@                        H�4H�4@z�5��(@y%jW�vH@H�4H�4@;��,��@;l��F:B@0#0#�?��#�� @                z�5��@<l��F:B@0#0#�?z�5��@��/���@0#0#�?        �cp>@        z�5��@��/����?0#0#�?z�5��@                        ��/����?0#0#�?        ��/����?                        0#0#�?        On��O@@        ���>��@��On�(@��+��+@z�5��@��On�(@0#0#�?;��,��@�cp>@0#0#�?                0#0#�?;��,��@�cp>@        ;��,��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#��@                        ��/����?        ��#���?0����/#@                D�JԮD!@        ��#���?��/����?                ��/����?        ��#���?                ��#���?        0#0#@                0#0#@��#���?                        ��/���@dJ�dJ�A@        �cp>@=�C=�C?@        ��/����?                ��/����?=�C=�C?@        ��/����?�;�;;@        ��/����?                        �;�;;@        ��/����?0#0#@                0#0#@        ��/����?                0����/@0#0#@                0#0#@        0����/@                0����/@                ��/����?                �cp>@        ��b:��:@�e�_��7@�z��z�R@�k(��2@E�JԮD1@eJ�dJ�A@��#��0@���-��*@H�4H�4@��#��0@���-��*@0#0#�?�P^Cy/@E�JԮD!@        �P^Cy/@0����/@        z�5��(@��/����?        ���>��@                ;��,��@��/����?                ��/����?        ;��,��@                z�5��@��/���@        ��#���?��/���@                ��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                        ��/���@        ��#���?0����/@0#0#�?        0����/@0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                �cp>@        ��#���?                                ��+��+@��#�� @��/���@�s?�s?=@        ��/���@�C=�C=<@        ��/���@H�4H�4(@        ��/����?                ��/����?H�4H�4(@                ��+��+$@        ��/����?0#0# @        ��/����?                        0#0# @                0#0#0@��#�� @        0#0#�?                0#0#�?��#�� @                ��#�� @���-��@������C@z�5��@                ��#�� @���-��@������C@        �cp>@0#0# @        �cp>@                        0#0# @��#�� @��/����?�z��z�B@��#�� @        H�4H�4@��#�� @                                H�4H�4@        ��/����?S2%S2%A@        ��/����?��+��+$@                ��+��+$@        ��/����?                        H�4H�48@��#���?��/����?��+��+$@��#���?��/����?                ��/����?        ��#���?                                ��+��+$@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��;hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK߅�h��B�0         r                 @@�?N�Ϭ;.�?&      ��pQ�}@       -                 Цx�?p,Z�J=�?�       0�#jl@       "                 �>fR?����S��?F       �a#6�[@                        P�<8?��.�?:       �2�x�PW@                        `xNv?�IF^ڰ�?.       �m���R@                          \��?X��e�)�?)       TVl��P@                         �JV�?��x_F-�?       y%jW�v8@                        ��V?�:�^���?       ��]�ڕ5@	                         ����?F���'0�?       �C�� T"@
                        "?`n����?       � ��w<@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �               z�5��@������������������������       �      �<       |�5��(@                        X��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?                        ��$?����N-�?       �#[�$E@������������������������       �        	       �P^Cy/@                        �Q�?h�s�	�?       g���:@                        ����?`n����?       � ��w<@������������������������       �               ��#�� @                         ���?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?                           �?      �<       <��,��4@������������������������       �               |�5��(@������������������������       �               ��#�� @                        pTF�?� �_rK�?       J�@��"@������������������������       �               ;��,��@������������������������       �      ��       ��/���@        !                 ����?*@ȱ��?       ���~1@������������������������       �      �<
       ��|��,@������������������������       �      ȼ       z�5��@#       ,                 �Us9?x �_rK�?       J�@��2@$       )                 @�eo?h��H��?
       v�I�+@%       &                  ��n?�`@s'��?       Ei_y,*@������������������������       �               ��/���@'       (                 ��,?b%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?*       +                 ����?�_�A�?       肵�e`@������������������������       �               ;��,��@������������������������       �      �<       ��/����?������������������������       �               ��#��@.       m                 ��ӱ?��Shޫ�?I       H�*�]@/       d                  ���?�lt��?B       e&��@Z@0       [                    �?<�e\�?6       ��K��T@1       T                   �x�?@����?#       ٭	���I@2       K                 PUҦ?��jT���?       ��6��E@3       >                 ��??�A�4qF�?       椫�u�>@4       5                 p��h?����W�?
       �`���@*@������������������������       �               z�5��@6       ;                 p���? �Z�ܙ�?       c����@7       :                 `�_{?�@G���?       hu��@8       9                 ݌��?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��/����?<       =                 `�ռ?Zn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @?       H                 ��J�?�v���?       mtL�	�1@@       G                 �5W�?��r�S�?       �f��%/@A       D                 �V"P?���k�L�?       sk��#@B       C                  `S��?      �<       ���-��@������������������������       �               ��/����?������������������������       �               0����/@E       F                  PV��?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?������������������������       �               �cp>@I       J                 �H��?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?L       M                  h��?�����?       �l�C�J)@������������������������       �               0#0# @N       S                 p���?�^�#΀�?       O�{��A%@O       P                 H�?ʔfm���?       ��Z�N@������������������������       �               ��#���?Q       R                 ���?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �      ��       ���-��@U       V                 ���?x^�(���?       � K�h @������������������������       �               ��#���?W       X                 hU�<?P�ih�<�?       ��
@������������������������       �               ��+��+@Y       Z                ��v�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?\       ]                 ��?J9�)\e�?       `���b@@������������������������       �               ��/���@^       _                 J�P?�����?       �O��8@������������������������       �               ��/����?`       c                 �{��?��v^�n�?       ��m�7@a       b                 p'v�?Zn����?       ~��Y-"@������������������������       �      ��       z�5��@������������������������       �               �cp>@������������������������       �      ��       ���>��,@e       f                 ����?
k�e���?       �	~�a5@������������������������       �               ��#�� @g       l                  [$�?�[nD���?
       ���y�O3@h       k                  0p��?Z%��̫�?       �@�o#@i       j                 p5W�?�;[��G�?       �O�;�]!@������������������������       �      �<       ��/���@������������������������       �               0#0#�?������������������������       �      ܼ       ��#���?������������������������       �               0����/#@n       q                   ҏ�?"���3�?       &��X&@o       p                 ���?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               0#0# @s       �                   �0�?�׉��s�?�       �yH㏼n@t       �                 `s5�?v���W�?N       ���	�&^@u       �                 ���?�*ӟC�?       ���$j�H@v       y                 �7/�?�L��;�?       mG�y;@w       x                 ��O�?jP�D�?       �A��P?$@������������������������       �      �<       ���>��@������������������������       �      ȼ       �cp>@z                         
�?�T`�[k�?       �m����0@{       ~                 @�?��E�B��?       dߞKC.@|       }                  ����?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0#@������������������������       �               vb'vb'"@������������������������       �      ȼ       ��/����?�       �                 h��1?����>�?       z6gZ
6@�       �                 ����?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 p?�?�?�0�!�?       a`�T�4@������������������������       �      ��	       0#0#0@�       �                 ��c?��G���?       ��%�|@������������������������       �               ��/����?�       �                  ��?|��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?�       �                   ҏ�?	�{���?2       7�g�k�Q@�       �                 �U��?xLU���?       i�ҹ^�@������������������������       �               ���-��@������������������������       �               0#0#�?�       �                 �]�?={��L��?-       �,�O@�       �                 ����?\om`m�?       �N�h�oB@�       �                 NK�X?�7���?       S��"Xk@@�       �                 ����?|��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?�       �                    �?�A�o�?       j����=@�       �                 ��C�?g�wy��?       �f0�v&@������������������������       �               ;��,��@�       �                 ����?�g�vw�?       �Aws}8@�       �                 `��?r�T���?       ��e[�&@�       �                 ˃��?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �               0#0# @������������������������       �      ��       �k(��2@������������������������       �               0#0#@�       �                 ���?��dn��?       ͚?]��:@�       �                 *�}?dV�\Ga�?
       q�6t%@������������������������       �               0#0# @�       �                    �?)���?       x��uk!@�       �                ��Sl�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       ���-��@�       �                 p��?�¿���?       Hb0�*0@�       �                 �{��?T����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @�       �                   s��?���MF�?       �`�I-*@�       �                 �-�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 ��޲?�,m:��?	       ܃���=&@������������������������       �               �C=�C=@�       �                 �@��?f,���O�?       ���/>@������������������������       �               0#0# @�       �                  �Ԧ�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?�       �                 ��?�t�V���?I       m�ɼ~R_@�       �                  ��a?d�����?       gCS,bG@�       �                 08Y�?k��A�?       �r��6@�       �                 x��?Hy��]0�?       ���y"@������������������������       �               0#0#@�       �                  `%+�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 pa��?d�Ѿ�?       ޓr�0@�       �                    �?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @�       �                 �`��?�;�a
=�?
       ��l��+@�       �                 �&6�?�+�z���?	       LGh��
)@������������������������       �               �cp>'@������������������������       �               0#0#�?������������������������       �               0#0#�?������������������������       �               H�4H�48@�       �                 0���?�k=$�?,       �Q�&x�S@�       �                 p'v�?0,�#6?�?#       Z��̿.N@������������������������       �               %S2%S27@�       �                 p��J?�c3Q�I�?       �p+:��B@������������������������       �               vb'vb'2@�       �                 �?�?*�
Fq�?       /��3@�       �                 �j��?�~�&��?       >�]��@������������������������       �               ��/����?�       �                 ���?�AP�9��?       i��6��@������������������������       �               H�4H�4@�       �                  p�Z?|�G���?       ��%�|@������������������������       �               ��/����?�       �                 8���?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               #0#0&@�       �                 �-�?�gV8c��?	       "� a(2@������������������������       �               ��#�� @�       �                 ��?r����?       Qz�i0@������������������������       �               ��/����?������������������������       �      ��       �A�A.@�t�b�     h�hhK ��h��R�(KK�KK��h �B�  �����c@�-����`@�P��f@�Gp�=]@�'�xr�V@��+��+4@������S@Qn��O@@        Gy�5Q@��On�8@        �P^CyMP@鰑%@        Lp�}N@���-��@        ������3@0����/@        ������3@��/����?        ���>��@��/����?        ��#��@��/����?        ��#��@                        ��/����?        z�5��@                |�5��(@                        �cp>@                ��/����?                ��/����?        ��k(/D@��/����?        �P^Cy/@                {�5��8@��/����?        ��#��@��/����?        ��#�� @                ��#�� @��/����?        ��#�� @                        ��/����?        <��,��4@                |�5��(@                ��#�� @                ;��,��@��/���@        ;��,��@                        ��/���@        z�5��@��|��,@                ��|��,@        z�5��@                <��,��$@��/���@        z�5��@��/���@        ��#���?�cp>@                ��/���@        ��#���?��/����?        ��#���?                        ��/����?        ;��,��@��/����?        ;��,��@                        ��/����?        ��#��@                f:��,&C@��|��L@��+��+4@�k(��B@�a#6�K@H�4H�4(@Fy�5A@3����/C@#0#0&@��b:��*@���-��:@#0#0&@{�5��(@�cp>�9@��+��+@[Lg1��&@On��O0@H�4H�4@��#�� @��/���@0#0#�?z�5��@                ��#�� @��/���@0#0#�?        �cp>@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?        ��#�� @��/����?                ��/����?        ��#�� @                z�5��@��On�(@0#0# @��#���?��On�(@0#0# @��#���?���-��@0#0# @        ���-��@                ��/����?                0����/@        ��#���?        0#0# @                0#0# @��#���?                        �cp>@        ��#�� @                ��#���?                ��#���?                ��#���?0����/#@0#0# @                0#0# @��#���?0����/#@        ��#���?�cp>@        ��#���?                        �cp>@                ��/����?                ��/����?                ���-��@        ��#���?��/����?H�4H�4@��#���?                        ��/����?H�4H�4@                ��+��+@        ��/����?0#0#�?        ��/����?                        0#0#�?<��,��4@�cp>'@                ��/���@        <��,��4@��/���@                ��/����?        ;��,��4@�cp>@        z�5��@�cp>@        z�5��@                        �cp>@        ���>��,@                z�5��@E�JԮD1@0#0#�?��#�� @                ��#���?E�JԮD1@0#0#�?��#���?��/���@0#0#�?        ��/���@0#0#�?        ��/���@                        0#0#�?��#���?                        0����/#@        ��#���?��/����?0#0# @��#���?��/����?        ��#���?                        ��/����?                        0#0# @<��,��D@h
��F@�|˷|d@�k(��B@���-��:@�C=�C=L@���>��@/����/#@0#0#@@���>��@���-��@��8��8*@���>��@�cp>@        ���>��@                        �cp>@                ��/���@��8��8*@        ��/����?��8��8*@        ��/����?0#0#@        ��/����?                        0#0#@                vb'vb'"@        ��/����?                �cp>@��)��)3@        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?vb'vb'2@                0#0#0@        ��/����?0#0# @        ��/����?                ��/����?0#0# @                0#0# @        ��/����?        Lp�}>@D�JԮD1@H�4H�48@        ���-��@0#0#�?        ���-��@                        0#0#�?Lp�}>@鰑%@%S2%S27@�#���9@��/����?vb'vb'"@�#���9@��/����?��+��+@        ��/����?0#0# @                0#0# @        ��/����?        �#���9@��/����?H�4H�4@���>��@��/����?H�4H�4@;��,��@                ��#�� @��/����?H�4H�4@��#�� @��/����?0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?��#�� @                                0#0# @�k(��2@                                0#0#@��#��@D�JԮD!@�C=�C=,@��#���?��/���@0#0# @                0#0# @��#���?��/���@        ��#���?��/����?                ��/����?        ��#���?                        ���-��@        z�5��@��/����?H�4H�4(@��#�� @        0#0#�?                0#0#�?��#�� @                ��#���?��/����?#0#0&@        ��/����?0#0#�?                0#0#�?        ��/����?        ��#���?        ��+��+$@                �C=�C=@��#���?        H�4H�4@                0#0# @��#���?        0#0#�?��#���?                                0#0#�?��#��@D�JԮD1@�Wx�W�Y@��#�� @���-��*@=�C=�C?@��#�� @���-��*@�C=�C=@        ��/����?��+��+@                0#0#@        ��/����?0#0#�?        ��/����?                        0#0#�?��#�� @��On�(@0#0# @��#�� @��/����?                ��/����?        ��#�� @                        �cp>'@0#0# @        �cp>'@0#0#�?        �cp>'@                        0#0#�?                0#0#�?                H�4H�48@��#�� @��/���@xb'vb'R@        �cp>@�[��[�L@                %S2%S27@        �cp>@T2%S2%A@                vb'vb'2@        �cp>@0#0#0@        �cp>@��+��+@        ��/����?                ��/����?��+��+@                H�4H�4@        ��/����?0#0# @        ��/����?                ��/����?0#0# @        ��/����?                        0#0# @                #0#0&@��#�� @��/����?�A�A.@��#�� @                        ��/����?�A�A.@        ��/����?                        �A�A.@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJS�)/hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKÅ�h��B�*         �                  b?�@���7�?%      �!s���}@       �                 @���?4��Js�?�       
Tm�Iv@       n                 ����?�B=���?�       (���Xt@       c                  ��?����b�?�       ����l@       L                 P^N<?�Lա��?�       ���-�,i@                        `��`?ŀY���?f       ʍg$��c@                         ,v�>.µ*A
�?       ��A抌9@������������������������       �               ;��,��@	                          .p�?�`@s'��?       �[�_4@
                        hf�?z�����?       �4^$4�#@������������������������       �               0����/@                        0�?ܗZ�	7�?       j~���@������������������������       �               z�5��@������������������������       �      �<       ��/����?                         �9��?      �<       鰑%@������������������������       �               ��/����?������������������������       �               0����/#@       C                 ~`����$% �?W       �O��W�`@                         �Q�?v�h��?7       |�|vQ�U@                       D䔶�?��3Fi�?       :�"Ξs@������������������������       �               ��#�� @������������������������       �               ��+��+@       6                 p_Q�?�|��$��?4       	ǚ��S@       5                 @��?�ĕ��?"       �`� cG@       "                  �_�?v`f����?!       ��]��`F@       !                  ����?�=vo�`�?       �M��Jg/@                        U��?rR����?       p\����!@                        `s5�?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?                         �\͵?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �      ��       ���-��@#       (                 ��cy?#qGN��?       6|�<=@$       %                 �j��?�FO���?       �ߌ$@������������������������       �      ��       z�5��@&       '                �3�q?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@)       0                  ��^�?�F�?!�?       3V���2@*       +                 �/t?���/��?	       @z$S��'@������������������������       �               z�5��@,       -                  �Q�?f%@�"�?       �6�E�!@������������������������       �               0����/@.       /                 4Ń?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@1       4                 pTF�?��[����?       Hl�_A@2       3                 8?��?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               ��/���@������������������������       �               0#0# @7       B                 ���?��M��?       X��%U@@8       9                  �.�?����P�?       j����>@������������������������       �               �cp>@:       ;                 8LSR?�/B����?       �;�7��;@������������������������       �               ��/����?<       ?                 �|��?�z;/2�?       �=�X��9@=       >                 �?      �<	       ���>��,@������������������������       �               ��#�� @������������������������       �               {�5��(@@       A                 @��x?l7Y���?       ���r�&@������������������������       �               0#0#�?������������������������       �               ;��,��$@������������������������       �               0#0# @D       I                 �u�?��DN�?        QW�1��G@E       H                 ���p? v+]�7�?       p�vc��D@F       G                 �G�o?X�j���?	       ���z"@������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?������������������������       �               ���b:@@J       K                 (v?      �<       �cp>@������������������������       �               ��/����?������������������������       �               0����/@M       \                 ���?������?       ��8%�E@N       W                    �?�Äy�?       ����B@O       P                  �Q�?h%@�"�?       ��[�7@������������������������       �               ��On�(@Q       V                  Pmj�?���Ѯ�?       ��GQ&@R       S                 h%B`?ʔfm���?       ��Z�N@������������������������       �               ��#���?T       U                 �ޥW?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �      �<       ���>��@X       [                 P��?@��c`�?	       %��t5)@Y       Z                 _��>f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �      ��       0����/#@]       b                 �5P?ģ���c�?       �>�!J!@^       a                 ��|?�zœ���?       IG���t@_       `                    �?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?d       g                 ��=�?�U����?       �b�:�7@e       f                p�<��?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?h       k                 0vb�? �����?       �ڬ�ڬ4@i       j                 02|+?T����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @l       m                 `��?      �<       ��,���1@������������������������       �               ��#���?������������������������       �               ��#��0@o       �                 ���?�S�m�!�?7       �܋[$Y@p       }                 �U�<?V& ��?       �WI�_I@q       r                 �~Ͱ?:�4�$�?       8�詬i7@������������������������       �               z�5��@s       t                   E(�?�x�nF}�?	       ��+#�N4@������������������������       �               ��#�� @u       v                 @N��?~��Z�{�?       i#��<2@������������������������       �               0#0# @w       z                 0���?�i^�c�?       �D9�V$@x       y                ��?��?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@{       |                 ����?�o���?       o�9�F@������������������������       �               0#0#@������������������������       �               ��#���?~       �                 �y�?d�t�v�?       �}���U;@       �                 �Q�?�����o�?       ^���v<3@������������������������       �               ��|��,@�       �                  �p�?���mf�?       毠�?b@������������������������       �      �<       ��/���@������������������������       �               0#0#�?�       �                 p���?�t����?       b�=�2 @������������������������       �               ��/����?�       �                  �^��?�.�KQu�?       �K̎@������������������������       �               z�5��@������������������������       �               0#0#@�       �                 �o�??<�����?       ��m{�H@�       �                  �Ѱ? LX�a��?       �����?@@�       �                 @*t3?�@G���?       hu��/@�       �                 (I��?���mf�?       �qB_-@�       �                    �?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               鰑%@������������������������       �               0#0#�?�       �                 ��N�?�=�z��?
       IS��0@������������������������       �               ��#�� @�       �                 ����?x��`p��?       T����-@�       �                 @ �?z�G���?       �֔�Э#@������������������������       �               �cp>@�       �                  �G?�?�AP�9��?       i��6��@������������������������       �               ��/����?������������������������       �               ��+��+@������������������������       �               ��+��+@�       �                 ��>�?1�~��?	       r��GQ1@������������������������       �               ��|��,@�       �                    �?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 PR��?L��fz�?       s�%�?@�       �                   �P�?�;�a
=�?       ��l��@������������������������       �               �cp>@�       �                  ����?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@�       �                  ���? a�ox��?       ���e�H8@�       �                p�~�?�J���?       a���@������������������������       �               0#0#�?�       �                 ���?�|2N��?       �3K}@������������������������       �               ��#�� @�       �                 �{��?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?������������������������       �               vb'vb'2@�       �                 `�0z?�v	����?E       �6����\@�       �                 ��f?tL�0���?       P~�)��2@������������������������       �               ��#���?�       �                  cy?d����?       �����1@�       �                 Ў m?�Jn�� �?       �+�i�0@�       �                 �<��?$^�yU�?       ��7�1�#@������������������������       �               ��+��+@�       �                 f?d�4���?       �tCP��@������������������������       �               0#0# @������������������������       �               �cp>@������������������������       �               �C=�C=@������������������������       �      �<       ��/����?�       �                  ��?@��
�?7        WJ;]1X@������������������������       �      ��       �s?�s?M@�       �                 �!�?�ދ��?       :UF#C@�       �                 0E��?d*�'=P�?        �2"@������������������������       �               0#0# @������������������������       �      ȼ       ��/����?�       �                 �)Ì?      �<       �s?�s?=@������������������������       �               0#0#�?������������������������       �               �C=�C=<@�t�bh�hhK ��h��R�(KK�KK��h �BH  ��Gp_b@U<�œb@�P��f@�5��P>b@M!��a@gJ�dJ�Q@������a@�-����`@H�4H�4H@Ky�5�_@��-��bT@0#0#0@��b:��Z@h
���S@�C=�C=,@�,����W@q��F:lI@��8��8*@��#�� @D�JԮD1@        ;��,��@                z�5��@D�JԮD1@        z�5��@���-��@                0����/@        z�5��@��/����?        z�5��@                        ��/����?                鰑%@                ��/����?                0����/#@        �k(���U@�-����@@��8��8*@����JG@���-��:@��8��8*@��#�� @        ��+��+@��#�� @                                ��+��+@�GpAF@���-��:@0#0# @������3@h
��6@��+��+@������3@h
��6@H�4H�4@��#��@鰑%@0#0#�?��#��@��/���@0#0#�?��#��@��/����?        ��#��@                        ��/����?                �cp>@0#0#�?        �cp>@                        0#0#�?        ���-��@        �P^Cy/@�cp>'@0#0# @�k(��"@��/����?        z�5��@                z�5��@��/����?                ��/����?        z�5��@                z�5��@鰑%@0#0# @z�5��@�cp>@        z�5��@                z�5��@�cp>@                0����/@        z�5��@��/����?                ��/����?        z�5��@                        0����/@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @        ��/���@                        0#0# @z�5��8@0����/@H�4H�4@{�5��8@0����/@0#0#�?        �cp>@        z�5��8@��/����?0#0#�?        ��/����?        z�5��8@        0#0#�?���>��,@                ��#�� @                {�5��(@                <��,��$@        0#0#�?                0#0#�?;��,��$@                                0#0# @��k(/D@���-��@        ��k(/D@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ���b:@@                        �cp>@                ��/����?                0����/@        z�5��(@��|��<@0#0#�?�k(��"@���-��:@        ��#�� @��/���.@                ��On�(@        ��#�� @�cp>@        ��#���?�cp>@        ��#���?                        �cp>@                ��/����?                ��/����?        ���>��@                ��#���?�cp>'@        ��#���?��/����?                ��/����?        ��#���?                        0����/#@        z�5��@��/����?0#0#�?z�5��@        0#0#�?��#���?        0#0#�?��#���?                                0#0#�?��#�� @                        ��/����?        ������3@��/����?0#0# @        ��/����?0#0#�?                0#0#�?        ��/����?        ������3@        0#0#�?��#�� @        0#0#�?                0#0#�?��#�� @                ��,���1@                ��#���?                ��#��0@                �P^Cy/@f#6�aJ@0#0#@@��b:��*@%jW�v%4@S2%S2%1@<��,��$@��/����?H�4H�4(@z�5��@                ���>��@��/����?H�4H�4(@��#�� @                ;��,��@��/����?H�4H�4(@                0#0# @;��,��@��/����?0#0#@��#��@��/����?                ��/����?        ��#��@                ��#���?        0#0#@                0#0#@��#���?                z�5��@/����/3@��+��+@        ;l��F:2@0#0#�?        ��|��,@                ��/���@0#0#�?        ��/���@                        0#0#�?z�5��@��/����?0#0#@        ��/����?        z�5��@        0#0#@z�5��@                                0#0#@��#�� @Qn��O@@�A�A.@��#�� @Nn��O0@�C=�C=,@        �cp>'@0#0#@        �cp>'@H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@        鰑%@                        0#0#�?��#�� @0����/@��+��+$@��#�� @                        0����/@��+��+$@        0����/@��+��+@        �cp>@                ��/����?��+��+@        ��/����?                        ��+��+@                ��+��+@        On��O0@0#0#�?        ��|��,@                ��/����?0#0#�?                0#0#�?        ��/����?        z�5��@�cp>@#0#06@        �cp>@0#0#�?        �cp>@                �cp>@0#0#�?                0#0#�?        �cp>@        z�5��@        ��-��-5@z�5��@        H�4H�4@                0#0#�?z�5��@        0#0# @��#�� @                ��#���?        0#0# @                0#0# @��#���?                                vb'vb'2@��#���?0����/@�����{[@��#���?��/���@�C=�C=,@��#���?                        ��/���@�C=�C=,@        �cp>@�C=�C=,@        �cp>@�C=�C=@                ��+��+@        �cp>@0#0# @                0#0# @        �cp>@                        �C=�C=@        ��/����?                ��/����?D�s?��W@                �s?�s?M@        ��/����?�z��z�B@        ��/����?0#0# @                0#0# @        ��/����?                        �s?�s?=@                0#0#�?                �C=�C=<@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ[س=hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK˅�h��Bh,         �                 0�0�?y�sy�T�?2      K�P&�}@       S                 @�(�?>x`3��?�       ����0�t@       "                 ��l?�2�.%�?{       �c�e�g@                        0��>]�Jm�?$       өhǫO@������������������������       �               E�JԮD!@       	                 `�]?X�	��`�?        ��U��J@                         �.�?\����?       P	K��@������������������������       �               ��/����?������������������������       �               z�5��@
                        ���r?n�)	C��?       T���/G@                        ��-�?���S�m�?       �[O�L�D@                        ���Q?�|2N��?       �3K}@������������������������       �               z�5��@������������������������       �               0#0# @                          B�?h���M�?       ���g�	B@                         խ�?�z�BC��?       �jϦ%�A@                        ���Y?L�gAW��?       �z��;@������������������������       �               鰑%@                        `&�k?>3#܅�?
       ���A�0@                        ��j�?���/��?       @z$S��@������������������������       �               �cp>@������������������������       �               z�5��@������������������������       �               鰑%@                        ���R?@��X�&�?       �6��	�@������������������������       �               �cp>@                         ���?�nɵ��?       Cad�J@������������������������       �               z�5��@                       @5	{�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      �<       ��#���?        !                  �.�?      �<       ;��,��@������������������������       �               ��#�� @������������������������       �               z�5��@#       R                 ��'�?�j�n�?W       �r\�u�_@$       I                 @F�D�0�=�?T       x*�m-^@%       8                 Цx�?�3I^���?A       Y�����V@&       5                  �tx?������?+       ���ѫO@'       0                 pM�D?�]���?&       �j0�W�L@(       /                 �94W?�����?#       +d�HI@)       .                 @�AV?DBms�?       ��֖��;@*       +                 �\И?`7uV��?        m}�'�:@������������������������       �               �,����7@,       -                 �R�־dn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               \Lg1��6@1       2                 `��?z��H��?       v�I�@������������������������       �               ��/����?3       4                 �Dph?��Z�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@6       7                  `s�?�@ȱ��?       nm���S@������������������������       �      ��       0����/@������������������������       �               ��#���?9       H                 ��=�?Vח���?       3��bXL<@:       A                    �?�)��R=�?       �
3�e19@;       @                  T?ܜ�x�?       e��إV3@<       =                   ��?�O
�*Q�?       �͉V�M2@������������������������       �               ��/���.@>       ?                 P��?h%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      �<       ��#���?B       C                 H�{�?�� ��?       qp� k@������������������������       �               �cp>@D       E                  ��?x��`p��?       �����@������������������������       �               0#0#�?F       G                  ��d�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ȼ       z�5��@J       O                 �7\?��=�Sο?       ����<@K       N                 x��?`7uV��?       m}�'�:@L       M                 �~�?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �               �k(���5@P       Q                 �uv?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      �       H�4H�4@T       a                 �!�?p��R��?[       3`���b@U       \                 ���?b����?       ��F{��:@V       W                 �N�~?�?�0�!�?
       a`�T�4@������������������������       �               ��/����?X       Y                 ���?8L�0�h�?	       k�e�3@������������������������       �      ��       ��8��8*@Z       [                    �?Hy��]0�?       ���y"@������������������������       �               ��+��+@������������������������       �      ȼ       ��/����?]       `                 pE	�?�w��d��?       �0���s@^       _                  ��?���mf�?       毠�?b@������������������������       �      �<       ��/���@������������������������       �               0#0#�?������������������������       �               0#0# @b       m                   .p�?0n��#�?M       C�Rp]@c       j                 �U��>�XӐ���?       ]�W=�3B@d       i                 `��?Xn����?       ��Y-2@e       h                 @tܣ?��k{��?	       _;�W� *@f       g                 P]ڒ?F���'0�?       �C�� T"@������������������������       �               ��/����?������������������������       �      ��       ���>��@������������������������       �      ȼ       ��/���@������������������������       �      Լ       ;��,��@k       l                    �?      �<       ;l��F:2@������������������������       �               0����/#@������������������������       �               E�JԮD!@n       �                 ���?��O���?6       
I4/VT@o       �                 �ve�?΄y&��?"       ��G��J@p       �                 @Z!�?\��$�?       �9a �E@q       r                   E(�?4���?       k�A@������������������������       �               ��#���?s       |                  ��~?�ص����?       ���O�A@t       {                 `Hx?�
�CX�?       ��:.�%@u       v                  P���?Ȕfm���?       ��Z�N@������������������������       �               �cp>@w       z                 �h�v?4=�%�?       �(J��@x       y                 �&%r?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      �<       ��/����?������������������������       �               H�4H�4@}       ~                    �?�F���?       ;�.�-7@������������������������       �               ��On�(@       �                 0��?V�ђ���?	       �oFݜh%@�       �                 3��?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ��       ��/���@�       �                 ����?r��`p��?       f;3@��!@������������������������       �               0#0#@�       �                 ��K�?l�4���?       �tCP��@������������������������       �               �cp>@������������������������       �               0#0# @�       �                 ��L�?\���'0�?       �C�� T"@������������������������       �               ���>��@������������������������       �      �<       ��/����?�       �                 �gY�?H���԰?       �����0<@������������������������       �      ��       �;�;;@������������������������       �      �<       ��/����?�       �                   ��?��^)&�?\       @���Ua@�       �                 `N�?��C��?D       ]O���X@�       �                  '�?X:}k�:�?        ��G@�       �                 x6v�?~���Y1�?       Fn���D@�       �                 ���6?t�GZ��?       O+A2?@�       �                 �#�?bn����?       ����45@������������������������       �        
       ��b:��*@�       �                    �?��r{��?       e�6� @������������������������       �               ��#���?������������������������       �               ���-��@�       �                 p�O�?X@ �F��?       tռ7�#@������������������������       �               H�4H�4@�       �                 P7&E?�`@s'��?       Ei_y,*@�       �                  H?��?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��/���@�       �                 ��vv?      �<       vb'vb'"@������������������������       �               0#0#�?������������������������       �               0#0# @�       �                 �Ô�?@y��]0�?       ���y"@������������������������       �               ��+��+@������������������������       �      ȼ       ��/����?�       �                 p�{�?Ʃwɰ��?$       ��	NȢJ@�       �                    �?��Y�?       �.	-21@�       �                 �}B�?T����1�?       ��;9�@������������������������       �               0#0# @������������������������       �               ��#��@�       �                 �oW�?�it�R��?	       ��ǿ%@������������������������       �               H�4H�4@�       �                  ����?���`�?       ��
�Me@������������������������       �               �cp>@�       �                 ����?��`i��?       �؛.�@������������������������       �               ��/����?�       �                  �!�?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?�       �                 �bW�?�/y߃�?       Va�7�B@�       �                  ���?��-}��?
       8�g51@�       �                 �j��?t�+(�s�?	       ��iq
6.@������������������������       �               ��+��+$@�       �                 `Z�?:�N9���?       ��{j�@�       �                 h�~�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               ��#���?������������������������       �      ȼ       ��/����?�       �                  =�a?�Qׅ؛�?       s�W)73@�       �                 ����?�J���?       ��*]Y@������������������������       �               ��#�� @������������������������       �               0#0# @������������������������       �      �<	       �A�A.@�       �                  H�?(����?       K�t@ħC@������������������������       �        
       ��)��)3@�       �                 @�/�?t�h�ku�?       �����%4@�       �                  ��?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?�       �                 ���?�#Vn\��?       I�~B�2@������������������������       �               ��/����?������������������������       �               S2%S2%1@�t�bh�hhK ��h��R�(KK�KK��h �B  ��b:��c@�JԮDmc@�|˷|d@�,���n`@����/�`@U2%S2%Q@z�YL�Z@����z�Q@#0#0&@�k(���5@�+Q��B@H�4H�4@        E�JԮD!@        �k(���5@��|��<@H�4H�4@z�5��@��/����?                ��/����?        z�5��@                �P^Cy/@�a#6�;@H�4H�4@<��,��$@�a#6�;@H�4H�4@z�5��@        0#0# @z�5��@                                0#0# @���>��@�a#6�;@0#0#�?z�5��@�a#6�;@0#0#�?z�5��@�e�_��7@                鰑%@        z�5��@���-��*@        z�5��@�cp>@                �cp>@        z�5��@                        鰑%@        z�5��@��/���@0#0#�?        �cp>@        z�5��@��/����?0#0#�?z�5��@                        ��/����?0#0#�?        ��/����?                        0#0#�?��#���?                ;��,��@                ��#�� @                z�5��@                ���#8U@�-����@@0#0# @���#8U@�-����@@0#0# @���>��L@�]�ڕ�?@0#0# @U^CyeJ@鰑%@        �#���I@�cp>@        5��tSH@��/����?        
�#���9@��/����?        
�#���9@��/����?        �,����7@                ��#�� @��/����?                ��/����?        ��#�� @                        ��/����?        \Lg1��6@                z�5��@��/���@                ��/����?        z�5��@��/����?                ��/����?        z�5��@                ��#���?0����/@                0����/@        ��#���?                ;��,��@鰑5@0#0# @��#�� @鰑5@0#0# @��#�� @E�JԮD1@        ��#���?E�JԮD1@                ��/���.@        ��#���?��/����?        ��#���?                        ��/����?        ��#���?                        ��/���@0#0# @        �cp>@                ��/����?0#0# @                0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?z�5��@                ��b:��:@��/����?        �#���9@��/����?        ��#��@��/����?        ��#��@                        ��/����?        �k(���5@                ��#���?��/����?        ��#���?                        ��/����?                        H�4H�4@|�5��8@4����-O@�[��[�L@        �cp>@��-��-5@        ��/����?vb'vb'2@        ��/����?                ��/����?vb'vb'2@                ��8��8*@        ��/����?��+��+@                ��+��+@        ��/����?                ��/���@H�4H�4@        ��/���@0#0#�?        ��/���@                        0#0#�?                0#0# @|�5��8@P!�ML@wb'vb'B@z�5��(@�e�_��7@        {�5��(@�cp>@        ���>��@�cp>@        ���>��@��/����?                ��/����?        ���>��@                        ��/���@        ;��,��@                        ;l��F:2@                0����/#@                E�JԮD!@        z�5��(@Pn��O@@vb'vb'B@z�5��(@�]�ڕ�?@vb'vb'"@;��,��@�_��e�=@vb'vb'"@;��,��@���-��:@H�4H�4@��#���?                ��#��@���-��:@H�4H�4@��#�� @�cp>@H�4H�4@��#�� @�cp>@                �cp>@        ��#�� @�cp>@        ��#�� @��/����?        ��#�� @                        ��/����?                ��/����?                        H�4H�4@��#�� @鰑5@                ��On�(@        ��#�� @E�JԮD!@        ��#�� @��/����?                ��/����?        ��#�� @                        ��/���@                �cp>@H�4H�4@                0#0#@        �cp>@0#0# @        �cp>@                        0#0# @���>��@��/����?        ���>��@                        ��/����?                ��/����?�;�;;@                �;�;;@        ��/����?        }�5��8@h
��6@ �q��V@�,����7@鰑5@�;�;K@�P^Cy/@���-��*@S2%S2%1@�P^Cy/@��On�(@H�4H�4(@�P^Cy/@��On�(@H�4H�4@���>��,@���-��@        ��b:��*@                ��#���?���-��@        ��#���?                        ���-��@        ��#���?�cp>@H�4H�4@                H�4H�4@��#���?�cp>@        ��#���?��/����?        ��#���?                        ��/����?                ��/���@                        vb'vb'"@                0#0#�?                0#0# @        ��/����?��+��+@                ��+��+@        ��/����?        ��#�� @��/���@�z��z�B@;��,��@0����/@�C=�C=@��#��@        0#0# @                0#0# @��#��@                ��#���?0����/@��+��+@                H�4H�4@��#���?0����/@0#0# @        �cp>@        ��#���?��/����?0#0# @        ��/����?        ��#���?        0#0# @                0#0# @��#���?                z�5��@�cp>@�A�A>@��#���?�cp>@��8��8*@��#���?��/����?��8��8*@                ��+��+$@��#���?��/����?H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@��#���?                        ��/����?        ��#�� @        S2%S2%1@��#�� @        0#0# @��#�� @                                0#0# @                �A�A.@��#���?��/����?�z��z�B@                ��)��)3@��#���?��/����?vb'vb'2@��#���?        0#0#�?��#���?                                0#0#�?        ��/����?S2%S2%1@        ��/����?                        S2%S2%1@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJnխphFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKͅ�h��B�,         �                 ��?)��T�?$      ��0(M~}@       {                 �"��?/��|�?�       �ru@       x                 �}]�?1��Km��?�       b���o@       k                  �/�?d]T�?�       �g��m@       P                 ���?�i�C8�?u       �ig�N�g@       1                 ���s?�@U�T�?]       �K��Xc@                        ��c?����q�?;       ��N0gW@                         �3��?̲�h�?        �+p |5@	       
                  �G?�?���/��?       U��7�@������������������������       �               ��/����?                        P�1?\n����?       � ��w<@������������������������       �               ��/����?                        ~`���d�$���?       �T�f@                         h��?bn����?       � ��w<@������������������������       �               ��#���?                        P�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#�� @                        0�2�?8e��}�?       ��Se+@������������������������       �      �<       �cp>'@                         `�J�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?       .                 �2OF?��h+�N�?+       ���20R@       +                 @R�v?�d�$���?&       �Cg�P@       (                 �kd1?@wE%h^�?"       ^�6m�1N@       !                 `.��>���d�0�?       Q8>�\E@                         P���?Zn����?       ~��Y-"@������������������������       �               ��/����?                         (u�?T����?       Q	K��@������������������������       �      �<       z�5��@������������������������       �      ȼ       ��/����?"       '                 �U���0�#�ݬ?       0X{Z�@@#       $                 ��V?h�j���?       ���z"@������������������������       �               ��/����?%       &                 ��Tv?      �<       ��#�� @������������������������       �               ��#��@������������������������       �               ��#��@������������������������       �               �,����7@)       *                 P��1?��{@��?       ��I�@2@������������������������       �               0����/@������������������������       �      ��       ��b:��*@,       -                 @�er?f%@�"�?       ��[�@������������������������       �      ��       ��/���@������������������������       �               ��#�� @/       0                 P>-l?8@ȱ��?       nm���S@������������������������       �      ��       0����/@������������������������       �               ��#���?2       M                 �C`�?��B�g��?"       ��絓�N@3       H                    �?rH����?        �쬥qJ@4       7                 J�e?"Q�aɴ�?       �Sy��A@5       6                   ҏ�?\����?       P	K��@������������������������       �               ��/����?������������������������       �               z�5��@8       =                   ���?TxO�gX�?       ����_<@9       <                  �\�?�3+�Pr�?
       Z-"�=L4@:       ;                 8�{?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               E�JԮD1@>       G                 ����?t�T���?       ��e[�& @?       D                 H?�26�
�?       5��*8E@@       A                   �x�?�d�$���?       �T�f@������������������������       �               ��#���?B       C                 �!�?����?       ��X�)B@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?E       F                 BQh�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               0#0#�?I       J                 �2FE?������?       �N0gX1@������������������������       �        	       ��|��,@K       L                  P�"�?j%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?N       O                 �#k�?      �<       ��#�� @������������������������       �               ��#��@������������������������       �               ��#��@Q       Z                  ��~�?�����?       �w�5G�B@R       S                  @V��?C�pB}��?       ����1$@������������������������       �               z�5��@T       U                  �g<�?���q���?       �:-ߩ�@������������������������       �               ��/����?V       Y                 ����?�nɵ��?       Cad�J@W       X                    �?����?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?������������������������       �               0#0#�?[       \                 �@�?`_"���?       ��hm�	;@������������������������       �               H�4H�4(@]       ^                 ����?��fܾ�?       z����-@������������������������       �               ��/����?_       f                    �?�n��T�?	       2~7�*@`       a                 X���?����]L�?       N66�ͯ@������������������������       �               ��#���?b       e                 �|�?�@G���?       hu��@c       d                 Lk�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               0#0#�?g       h                 `TԺ?a�ox��?       
c��0 @������������������������       �               ��#���?i       j                 �ڡs?      �<       �C=�C=@������������������������       �               0#0# @������������������������       �               ��+��+@l       w                 ���?�G|:=*�?       �`���G@m       t                 �SR�?t�j���?       �HI�G@n       q                 NK�X?��?	       ��l}�'*@o       p                  pjS�?d%@�"�?       ��[�@������������������������       �      ��       ��/���@������������������������       �               ��#�� @r       s                 0Ȳ�?d����?       P	K��@������������������������       �               ��/����?������������������������       �               z�5��@u       v                 ��F�?      �<       ��#��@@������������������������       �               ��#�� @������������������������       �               �P^Cy?@������������������������       �     ��<       0#0#�?y       z                   ҏ�?�*�'=P�?        �2"@������������������������       �               ��/����?������������������������       �               0#0# @|       �                 `�0z?�0��n�?;       ��O�pRV@}       ~                  ��{�?�y���@�?/       r;18�LR@������������������������       �               ��/���@       �                  8��?��h���?)       �=~Y�aP@�       �                 �b'�?>�VS�?'       p�M�PFO@�       �                   ҏ�?�{Bo(�?        �4�߬�I@������������������������       �               0#0#�?�       �                 �͡?Ҝf�&��?       �UΔKI@�       �                 ���?(�Zh�=�?       �"<2�C@�       �                 �Rˡ?4*V>��?       -�6B�@@�       �                 '4�h?ģ���c�?       �>�!J!@�       �                  @V��?��Z�	7�?       j~���@������������������������       �               z�5��@������������������������       �      �<       ��/����?������������������������       �               0#0#�?�       �                  �P�?pp!����?       �t��1�;@�       �                 H?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?�       �                 ��}?(�v���?       )f�n8@������������������������       �               0#0#�?������������������������       �               �cp>7@�       �                  �9��?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �               �cp>'@�       �                 ��?j�B��#�?       J[���%@�       �                 ����?�D�-,�?       �D'ŰO@������������������������       �               ��+��+@������������������������       �               ��#���?�       �                 Ђ��?& k�Lj�?       �q��l}@������������������������       �      ��       ��/���@������������������������       �               ��#���?�       �                 Tf��?P��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?�       �                 �Qï? s����?       Qz�i0@������������������������       �      ��
       ��8��8*@�       �                 ��!�?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                  @(B�?:�R߾�?R       �]2l��`@�       �                 `TF�?������?
       ���]�'@�       �                 p��?jQ��?       �s�=�!@������������������������       �      ��       �cp>@�       �                 �◓?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               H�4H�4@�       �                 ���?Pʪ'3��?H       P	'�^@������������������������       �               ;��,��@�       �                 `�4x?��*H�?G       �pX��]]@�       �                 pdJ�?4�Q$��?'       ��;�jAP@�       �                  @���?<�Xn��?       /MDD@�       �                 �fQ?�n���k�?       �-]ƗC@�       �                  uݝ?      �<       0#0#@@������������������������       �               0#0#�?������������������������       �               =�C=�C?@�       �                ���(z? �Qk��?       ��Th!�@�       �                 �$I�?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �               H�4H�4@������������������������       �      �<       ��#���?�       �                 ����?T�	j!�?       ��U�#�8@������������������������       �               ��/����?�       �                 0Ϯ�?$�����?        ۢ���6@������������������������       �               z�5��@�       �                 �x�L?lutee�?       P9��3@�       �                 ���?�@����?       ���a�#@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 @J�?d�4���?       �tCP��#@������������������������       �               0����/@�       �                 ��k�?�@����?       ���a�@�       �                 w?|��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �      ��       0#0# @�       �                 �+�[?      �<        ��8��8J@������������������������       �               0#0# @������������������������       �               #0#0F@�t�bh�hhK ��h��R�(KK�KK��h �B8  g:��,&c@������c@��+��+d@��tӹa@D�JԮDa@�[��[�L@�,���n`@鰑U@0#0#@@�,���n`@^�ڕ��T@H�4H�48@:��P^�V@������S@%S2%S27@�YLgqT@����z�Q@0#0# @Np�}N@�-����@@        ;��,��@On��O0@        ��#��@��/���@                ��/����?        ��#��@��/����?                ��/����?        ��#��@��/����?        ��#�� @��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                ��#�� @                ��#���?��On�(@                �cp>'@        ��#���?��/����?                ��/����?        ��#���?                �>��nK@E�JԮD1@        ��b:��J@��On�(@        �#���I@E�JԮD!@        e:��,&C@��/���@        z�5��@�cp>@                ��/����?        z�5��@��/����?        z�5��@                        ��/����?        ���b:@@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ��#��@                ��#��@                �,����7@                ��b:��*@0����/@                0����/@        ��b:��*@                ��#�� @��/���@                ��/���@        ��#�� @                ��#���?0����/@                0����/@        ��#���?                �k(���5@�+Q��B@0#0# @��b:��*@�+Q��B@0#0# @z�5��(@鰑5@0#0# @z�5��@��/����?                ��/����?        z�5��@                z�5��@&jW�v%4@0#0# @��#�� @;l��F:2@        ��#�� @��/����?                ��/����?        ��#�� @                        E�JԮD1@        ��#��@��/����?0#0# @��#��@��/����?0#0#�?��#��@��/����?        ��#���?                z�5��@��/����?        z�5��@                        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?                0#0#�?��#���?On��O0@                ��|��,@        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                ��#��@                ��#��@                ��#�� @��/���@��-��-5@z�5��@�cp>@0#0#�?z�5��@                z�5��@�cp>@0#0#�?        ��/����?        z�5��@��/����?0#0#�?z�5��@��/����?        z�5��@                        ��/����?                        0#0#�?��#�� @0����/@��+��+4@                H�4H�4(@��#�� @0����/@0#0# @        ��/����?        ��#�� @�cp>@0#0# @��#���?�cp>@0#0#�?��#���?                        �cp>@0#0#�?        �cp>@                ��/����?                ��/����?                        0#0#�?��#���?        �C=�C=@��#���?                                �C=�C=@                0#0# @                ��+��+@<��,��D@0����/@0#0#�?=��,��D@0����/@        ��#�� @0����/@        ��#�� @��/���@                ��/���@        ��#�� @                z�5��@��/����?                ��/����?        z�5��@                ��#��@@                ��#�� @                �P^Cy?@                                0#0#�?        ��/����?0#0# @        ��/����?                        0#0# @<��,��$@���-��J@k�6k�69@<��,��$@g#6�aJ@��+��+$@        ��/���@        ;��,��$@�'�xr�F@��+��+$@;��,��$@h
��F@0#0# @��#�� @'jW�v%D@H�4H�4@                0#0#�?��#�� @(jW�v%D@0#0# @��#�� @��|��<@0#0# @��#��@�a#6�;@0#0# @z�5��@��/����?0#0#�?z�5��@��/����?        z�5��@                        ��/����?                        0#0#�?��#���?�cp>�9@0#0#�?��#���?�cp>@                �cp>@        ��#���?                        �cp>7@0#0#�?                0#0#�?        �cp>7@        ��#��@��/����?                ��/����?        ��#��@                        �cp>'@        ��#�� @��/���@��+��+@��#���?        ��+��+@                ��+��+@��#���?                ��#���?��/���@                ��/���@        ��#���?                        ��/����?0#0# @                0#0# @        ��/����?                ��/����?�A�A.@                ��8��8*@        ��/����?0#0# @        ��/����?                        0#0# @\Lg1��&@1����/3@�Wx�W�Y@��#�� @���-��@H�4H�4@��#�� @���-��@                �cp>@        ��#�� @��/����?                ��/����?        ��#�� @                                H�4H�4@�k(��"@��On�(@n�6k�6Y@;��,��@                ��#��@��On�(@n�6k�6Y@��#��@��On�(@K�4H�4H@��#���?�cp>@wb'vb'B@        �cp>@xb'vb'B@                0#0#@@                0#0#�?                =�C=�C?@        �cp>@0#0#@        �cp>@0#0#�?        �cp>@                        0#0#�?                H�4H�4@��#���?                z�5��@/����/#@H�4H�4(@        ��/����?        z�5��@��/���@H�4H�4(@z�5��@                        ��/���@H�4H�4(@        ��/����?0#0# @        ��/����?                        0#0# @        �cp>@0#0#@        0����/@                ��/����?0#0#@        ��/����?0#0# @                0#0# @        ��/����?                        0#0# @                ��8��8J@                0#0# @                #0#0F@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�[�.hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKۅ�h��B�/         �                  ��?���tF?�?.      �b0c�}@       c                 ��H?t�]i�?�       '%1aC�q@       L                  ����?(����?       �����j@                        pt"?d `+��?Z       ���SBc@                         V�7?
KE��?       �-`R�B@                        x��?f����?       :��18>@                          \��?��h!��?       W�v%jW;@       	                 ,*������/��?	       K9U6�+@������������������������       �               0����/@
                        ��Yg?F���'0�?       �C�� T"@������������������������       �               ��/����?                           �?      �<       ���>��@������������������������       �               ��#���?������������������������       �               z�5��@                        �yW?l�s�	�?       e���*@������������������������       �               ��/����?������������������������       �               {�5��(@                        �sM?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?                        8*��?��|��?       ���ĺw@������������������������       �               ��#�� @������������������������       �      ��       0����/@       #                   ҏ�?������?D       m9O?]@       "                  ���?� �_rK�?       J�@��2@                        ��H�?d%@�"�?	       ��[�'@                        �m�?�`@s'��?       Ei_y,*@������������������������       �               ��/���@                         �0��?d%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?        !                 ��{?ܗZ�	7�?       j~���@������������������������       �               z�5��@������������������������       �      �<       ��/����?������������������������       �               z�5��@$       %                  9�>������?8       
�yz�X@������������������������       �               �cp>@&       K                 (�V�?4�|gv��?7       ��{�HX@'       ,                 �n5]?�4׼?��?6       �^�}��W@(       )                  �a�?f%@�"�?       ��[�@������������������������       �               �cp>@*       +                    �?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?-       4                 `�y�? Yjǯ�?2       �oBͦJV@.       /                 ��?����Y�?       3K}@�D@������������������������       �      ��       ��#��@@0       3                    �?��t1u�?       "�te!� @1       2                 Н�?T����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �      ��       ;��,��@5       H                 ��0�?�P��=�?       /�9�G@6       7                 �5W�?Z�]v\{�?       f�+'�D>@������������������������       �               ��#�� @8       C                  ��?�y��B�?       ��4��5@9       @                  `��? [��.��?       -���d.@:       =                 NK�X?vp�?�r�?       �E��
$@;       <                  �9��?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@>       ?                  �\~?�����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?A       B                 @�?      �<       ;��,��@������������������������       �               ��#�� @������������������������       �               z�5��@D       G                 P%W�?�`@s'��?       Ei_y,*@E       F                   ��?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��/���@I       J                 p\�?��:V��?
       �GP�1@������������������������       �        	       ��#��0@������������������������       �      �<       ��/����?������������������������       �     ��<       0#0#�?M       `                 ��G�?\���v�?%       dߟ���M@N       _                 �'U�?�W�W��?        �Zc���H@O       ^                 ��?"ذD���?       ������F@P       Y                 �]t?b�T��?       ��	�}FC@Q       V                 �y���rF9i5�?       l�HhH9@R       U                 �3�_?ʔfm���?       �0��z'@S       T                  ��?      �<       D�JԮD!@������������������������       �               ��/���@������������������������       �               0����/@������������������������       �      ȼ       z�5��@W       X                 ���@?�(߫$��?
       2H����*@������������������������       �               \Lg1��&@������������������������       �      ȼ       ��/����?Z       [                 �{k�?$e��}�?       ��Se+@������������������������       �      �<       鰑%@\       ]                 ����?^%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �               ���>��@������������������������       �               ��#��@a       b                  ��~?����h�?       @��o{#@������������������������       �               H�4H�4@������������������������       �      ��       ���-��@d       k                 ��,P?^��pqp�?,       �Tu��Q@e       h                 ��j�?�n�l���?       ���5F'@f       g                 p��?�;[��G�?       �O�;�]!@������������������������       �      �<       ��/���@������������������������       �               0#0#�?i       j                 �-�?V%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?l       }                  ��`?���C��?%       F��+~8M@m       |                 @F���_~"��?       ���Oo>@@n       o                 ����?���G���?       ]]���X<@������������������������       �               �cp>'@p       q                 �?b�o~��?
       �if^��0@������������������������       �               z�5��@r       y                 �y�?�Y�Z�?	       V�S��u+@s       t                  �<�?Δfm���?       ��Z�N@������������������������       �               �cp>@u       x                  �6��?
4=�%�?       �(J��@v       w                 �d"�?bn����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      �<       ��/����?z       {                 �V"P?x�G���?       '5L�`�@������������������������       �               �cp>@������������������������       �               H�4H�4@������������������������       �      ��       ��#��@~       �                 0��?ƎA���?       �l���9@       �                 ���?��íxq�?       $2��-�@�       �                  4#�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �      ��       ��/���@�       �                    �?�?�0�!�?       a`�T�4@������������������������       �      ȼ       �C=�C=,@�       �                 n~?���`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0#@�       �                   E(�?��K/���?�       �{�~�g@�       �                 �	�?��I<��?       Z���5�B@�       �                 �0��?���.�2�?       ��k	j3@�       �                 p���?j��H��?       v�I�@������������������������       �      ��       ��/���@������������������������       �               z�5��@�       �                 ��׍?      �<       ��On�(@������������������������       �               �cp>@������������������������       �               0����/#@�       �                 (=��?X�b���?
       �^Pb
2@�       �                 �!'�?@
:����?       {��"�%@�       �                 ��{�?��n��?       �-H�\@������������������������       �               ��/���@�       �                 @2��?��q�R�?       C}Ԥ@�       �                  ����?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �               ��#��@������������������������       �               �C=�C=@�       �                 pg_�?x�qm/A�?l       �M����b@�       �                 p��y?���)+��?X       N��#8�]@�       �                 GW�d?�:o��x�?6       ���R@�       �                 �j%?�ZX���?       QI�|�?@�       �                 ����?�x:o��?       r��L- 4@�       �                  ��u�?p�1���?       hD�LzF*@������������������������       �        
       H�4H�4(@������������������������       �      �<       ��#���?�       �                    �?�w��d��?       �0���s@������������������������       �               ��/����?�       �                 x�e�?~�G���?       '5L�`�@������������������������       �               �cp>@������������������������       �               H�4H�4@�       �                 �Q�?�֪u�_�?       ��?�8'@�       �                 p�)�?�}	;	�?       uK�>4%@������������������������       �               0����/#@������������������������       �               0#0#�?������������������������       �               0#0#�?�       �                  p��?\o�i�?       �s��mD@�       �                 ����?��,���?       \+ͮ�B@�       �                 ��?}��j�?       r$��Y5@�       �                 �]�?\�L�R��?       ��z��.@������������������������       �               ��/����?�       �                 `s5�?�b���:�?       �
#���,@�       �                 h��1?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      ��       [Lg1��&@�       �                 @� ?��]ۀ��?       E���O@������������������������       �               ��#���?�       �                 �mf�?�@����?       ���a�@������������������������       �               ��/����?������������������������       �               0#0#@�       �                    �?�p���K�?       C2(ߪ{0@�       �                  ��^�?D��NV=�?       �t�ܲ@�       �                 ��I�?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 �w��?�+�z���?       LGh��
)@������������������������       �               ���-��@�       �                 ���?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �               0����/@������������������������       �      �       H�4H�4@�       �                    �?|9��{�?"       �b�:�G@������������������������       �               ��-��-5@�       �                 8�C�?�N�+�?       ����:@�       �                  �Ԧ�?0�r��-�?       ���w�5@������������������������       �        	       H�4H�4(@�       �                  ��^�?d����?       �����!@������������������������       �               ��/����?������������������������       �      ��       �C=�C=@�       �                 f�?vutee�?       Q9��@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?�       �                 �M�?p=W�d��?       �q�գ*?@�       �                 p�?lutee�?       Q9��@�       �                 8��?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0# @������������������������       �               ��8��8:@�t�b�T     h�hhK ��h��R�(KK�KK��h �B�  ����bze@�B�)Dd@]x�WxEa@�k(��b@^#6�aZ@�s?�s?=@YUUUU5a@M!��Q@H�4H�4@
��G�[@'jW�v%D@H�4H�4@�k(���5@��/���.@        ������3@鰑%@        ������3@��/���@        ���>��@���-��@                0����/@        ���>��@��/����?                ��/����?        ���>��@                ��#���?                z�5��@                z�5��(@��/����?                ��/����?        {�5��(@                        �cp>@                ��/����?                ��/����?        ��#�� @0����/@        ��#�� @                        0����/@        �GpAV@��On�8@H�4H�4@;��,��$@��/���@        ��#��@��/���@        ��#���?�cp>@                ��/���@        ��#���?��/����?        ��#���?                        ��/����?        z�5��@��/����?        z�5��@                        ��/����?        z�5��@                ������S@E�JԮD1@H�4H�4@        �cp>@        ������S@��|��,@H�4H�4@������S@��|��,@0#0# @��#�� @��/���@                �cp>@        ��#�� @��/����?        ��#�� @                        ��/����?        f:��,&S@鰑%@0#0# @��k(/D@        0#0#�?��#��@@                ���>��@        0#0#�?��#�� @        0#0#�?                0#0#�?��#�� @                ;��,��@                �YLg1B@鰑%@0#0#�?������3@0����/#@0#0#�?��#�� @                \Lg1��&@0����/#@0#0#�?<��,��$@��/���@0#0#�?;��,��@��/���@0#0#�?        �cp>@0#0#�?                0#0#�?        �cp>@        ;��,��@��/����?        ;��,��@                        ��/����?        ;��,��@                ��#�� @                z�5��@                ��#���?�cp>@        ��#���?��/����?        ��#���?                        ��/����?                ��/���@        ��#��0@��/����?        ��#��0@                        ��/����?                        0#0#�?��b:��:@�_��e�=@H�4H�4@��b:��:@�cp>7@        \Lg1��6@�cp>7@        �P^Cy/@�cp>7@        ���>��,@鰑%@        z�5��@D�JԮD!@                D�JԮD!@                ��/���@                0����/@        z�5��@                \Lg1��&@��/����?        \Lg1��&@                        ��/����?        ��#���?��On�(@                鰑%@        ��#���?��/����?                ��/����?        ��#���?                ���>��@                ��#��@                        ���-��@H�4H�4@                H�4H�4@        ���-��@        ZLg1��&@����z�A@%S2%S27@��#���?0����/#@0#0#�?        ��/���@0#0#�?        ��/���@                        0#0#�?��#���?��/����?        ��#���?                        ��/����?        ;��,��$@�cp>�9@#0#06@�k(��"@%jW�v%4@H�4H�4@;��,��@%jW�v%4@H�4H�4@        �cp>'@        ;��,��@D�JԮD!@H�4H�4@z�5��@                ��#�� @D�JԮD!@H�4H�4@��#�� @�cp>@                �cp>@        ��#�� @�cp>@        ��#�� @��/����?        ��#�� @                        ��/����?                ��/����?                �cp>@H�4H�4@        �cp>@                        H�4H�4@��#��@                ��#���?�cp>@��)��)3@��#���?��/���@0#0#�?��#���?        0#0#�?��#���?                                0#0#�?        ��/���@                ��/����?vb'vb'2@                �C=�C=,@        ��/����?0#0#@        ��/����?                        0#0#@\Lg1��6@P!�ML@�;�;[@��#�� @鰑5@0#0# @z�5��@Nn��O0@        z�5��@��/���@                ��/���@        z�5��@                        ��On�(@                �cp>@                0����/#@        ;��,��@0����/@0#0# @;��,��@0����/@0#0#�?��#���?0����/@0#0#�?        ��/���@        ��#���?��/����?0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?        ��#���?                ��#��@                                �C=�C=@���>��,@����z�A@p�6k�6Y@���>��,@�-����@@p�fm��Q@���>��,@�_��e�=@�C=�C=<@��#���?���-��*@S2%S2%1@��#���?��/���@�A�A.@��#���?        H�4H�4(@                H�4H�4(@��#���?                        ��/���@H�4H�4@        ��/����?                �cp>@H�4H�4@        �cp>@                        H�4H�4@        /����/#@0#0# @        /����/#@0#0#�?        0����/#@                        0#0#�?                0#0#�?��b:��*@On��O0@#0#0&@��b:��*@On��O0@0#0# @z�5��(@�cp>@H�4H�4@[Lg1��&@��/����?0#0# @        ��/����?        \Lg1��&@��/����?0#0# @        ��/����?0#0# @        ��/����?                        0#0# @[Lg1��&@                ��#���?��/����?0#0#@��#���?                        ��/����?0#0#@        ��/����?                        0#0#@��#���?���-��*@0#0# @��#���?��/����?0#0#�?��#���?        0#0#�?                0#0#�?��#���?                        ��/����?                �cp>'@0#0#�?        ���-��@                0����/@0#0#�?                0#0#�?        0����/@                        H�4H�4@        ��/���@�
��
�E@                ��-��-5@        ��/���@#0#06@        ��/����?��)��)3@                H�4H�4(@        ��/����?�C=�C=@        ��/����?                        �C=�C=@        ��/����?H�4H�4@                H�4H�4@        ��/����?                ��/����?�s?�s?=@        ��/����?H�4H�4@        ��/����?0#0#�?                0#0#�?        ��/����?                        0#0# @                ��8��8:@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��=hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKh��BH4         �                 �H�?�0�*T�?(      ZX��؄}@       {                   �x�?�JOa�?�       ��$F5u@       X                 ����?E��ɵ��?�       �c��Bml@       ?                 ��??�W>�?p       9R���cg@       >                 �X��?d��/|��?T       �1�~ea@                         ��^�?x{|��?M       V	&���^@                        ��
?h�r{��?       e�6� @������������������������       �               0����/@	       
                  Pmj�?b%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?       =                 `=��?T�"L$#�?G       ��Ґ�\@                        �$?Z?@�G�1�?A       ��[Z@                        0�?& k�Lj�?	       e*�}#<-@                        �U�?Dǵ3���?       �q�ͨ�@                         �.�?ޗZ�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@������������������������       �      ��       �cp>@������������������������       �               ���-��@                          Mt?R�]v\{�?8       N�`���V@                        p�k?�v^�n�?       ��m�G@                         =�m?���+@�?       ���
$F@                        �6�b?���Ѯ�?       ��GQ&@������������������������       �               ��#�� @������������������������       �      ȼ       �cp>@                        @F�      �<       ��#��@@������������������������       �               Jp�}>@������������������������       �               z�5��@������������������������       �      �       �cp>@       :                  ���?nB�4|��?       ��?��E@        1                 NK�X?)���?       .zL<C@!       ,                  �JV�?�Ӏ�j�?       �~�5�d9@"       '                 P"ƭ?��b�}�?       ���\�#@#       &                    �?�d�$���?       �T�f@$       %                 �㚡?bn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               ��#�� @(       +                 @��?h�4���?       �tCP��@)       *                  ;�?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �               0#0#�?-       .                 �Ȕ�?����VV�?	       A�R.�.@������������������������       �               ��On�(@/       0                 �m�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?2       3                  �?��?	       ��l}�'*@������������������������       �               z�5��@4       5                  @mj�?��|��?       ���ĺw@������������������������       �               ��/���@6       7                  P���?^n����?       � ��w<@������������������������       �               ��#���?8       9                %I���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?;       <                 �MR�?      �<       ;��,��@������������������������       �               ��#���?������������������������       �               ��#��@������������������������       �               <��,��$@������������������������       �               ��b:��*@@       U                 .1�?������?       ���c�I@A       L                 @F�"~_h`�?       �d��F@B       I                  nl?ܜ�x�?       �-��=@C       H                 ���d?�O-r��?       �.w��e)@D       E                 x�S?�^�#΀�?       O�{��A%@������������������������       �               ��/���@F       G                 �.�\?\%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#�� @J       K                 ���@?      �<       On��O0@������������������������       �               E�JԮD!@������������������������       �               ��/���@M       R                 `��^?RR9�� �?	       ���55 0@N       O                 �U�K?ʔfm���?       ��Z�N@������������������������       �               ��#�� @P       Q                 �GE?      �<       �cp>@������������������������       �               �cp>@������������������������       �               �cp>@S       T                 ���~?�J���?       ��*]Y @������������������������       �               ��#��@������������������������       �               0#0#@V       W                 p_��?��|2N��?       �3K}@������������������������       �               z�5��@������������������������       �               0#0# @Y       b                   E(�?TOF�$�?       �E�ϴ&D@Z       a                 �=��?:4|���?       	�T|qt2@[       `                 �¼�?)���?       y��uk1@\       _                 ��?��i�@M�?       ���wzb0@]       ^                 �Q�?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �        	       ���-��*@������������������������       �      �<       ��#���?������������������������       �      �<       ��#���?c       p                  ��?cH-����?       q�c#��5@d       k                  ����?����h�?       @��o{#@e       j                ��ǳq?�;�a
=�?       ��l��@f       g                 py��?�@G���?       hu��@������������������������       �               ��/����?h       i                  L��?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               �cp>@l       m                ��X�p?z��`p��?       �����@������������������������       �               0#0#�?n       o                 PFe�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?q       x                 �
׭?�Z'Q���?       ���]�6(@r       s                 ����?�N̸��?       �#�zY9$@������������������������       �               H�4H�4@t       u                 ���?f,���O�?       ���/>@������������������������       �               0#0# @v       w                  �P��?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?y       z                 0�I�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?|       �                 �G�?��[{X��?F       l'P�Ob[@}       �                 ����?!�T��?0       �sك�S@~       �                 h�/s?� �c�?,       ų��(Q@       �                 0-3�?Z���L�?#       	گ�L@�       �                 ���@?��mS�w�?       ��@C@�       �                    �?\����?       R	K��<@�       �                 �@�?X\Cl[��?       >�s�d�9@�       �                  �d%�?xb8�Y�?       GJͰ8@�       �                  ���?pN:�*ط?       I�G�3@�       �                 �/��?|���X��?	       &��֞&@�       �                 ���>���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ��       �k(��"@������������������������       �               ��#�� @�       �                 �x�?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �      �<       ��/����?�       �                  �G?�?dn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @�       �                 0�2�?������?       �4^$4�#@�       �                 h��?      �<       ���-��@������������������������       �               ��/����?������������������������       �               �cp>@������������������������       �               z�5��@�       �                 �|T?�Jcү��?
       W��,3@�       �                 �4�X?7�H���?	       ǯ��02@������������������������       �               �cp>@�       �                 �S��?��2(&�?       �e4��\.@������������������������       �               �C=�C=@�       �                 X�P�?b,���O�?       ���/> @�       �                  ��^�?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?������������������������       �               ��+��+@������������������������       �      �<       ��#���?�       �                 P�J�?�^�F�M�?	       ��ޚ�&@������������������������       �               ��/����?������������������������       �               ��+��+$@�       �                  �Mm�?��fm���?       ��Z�N@�       �                    �?���/��?       V��7�@�       �                 (p�:?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      �<       ��/����?������������������������       �               ��/���@�       �                 Ȋ�8?Gb�����?       4g���@@�       �                 �#��?�_�A�?       炵�e`@�       �                    �?�����?       �O��@������������������������       �               ��#���?�       �                 ���?�d�$���?       �T�f@�       �                 ��R�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               z�5��@������������������������       �      ȼ       ��/����?�       �                  ���?�g���E�?       �m���9@�       �                 ����?z�G���?       �֔�Э#@�       �                 ���?�֪u�_�?       ��?�8@������������������������       �               �cp>@�       �                  �E�?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �               0#0#@������������������������       �        
       0#0#0@�       �                 `�4x?ܼ��=0�?U       q9)=G�`@�       �                 �;�?j)��T^�?3       uu��yT@�       �                 05D�?z2R}�-�?*       }(�D0P@�       �                 �4�?(l����?       �֕;Nu3@�       �                 �bl?.�(��?
       ��V-�*@�       �                ���E�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?�       �                 � 	�?|���X��?       '��֞&@������������������������       �               ��/����?������������������������       �      �<       ;��,��$@�       �                  z��?�D#���?       �B�j@������������������������       �               0#0#@������������������������       �               ��#�� @�       �                 h��?���k���?       e��F@�       �                 ��?Ի�$�+�?       u��;k4@�       �                  h��?�Qk��?       ��Th!�@������������������������       �               ��/����?�       �                 �n�b?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?�       �                    �?e��}�?       ��Se+@�       �                  P�"�?& k�Lj�?       �q��l}@�       �                 ����?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 �I�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               E�JԮD!@�       �                 �!ܳ?��lk��?       �:;��8@������������������������       �               ��+��+@�       �                 ����?N���|�?       �I0h��3@�       �                 ���?�T�"��?       ��`2�Z+@�       �                    �?�AP�9��?       i��6��@������������������������       �               0#0#@�       �                   �0�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �      ȼ       ���-��@�       �                 �\��?T����1�?       ��;9�@�       �                 ���?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               z�5��@�       �                 `
��?      �<	       S2%S2%1@������������������������       �               H�4H�4@������������������������       �               �C=�C=,@������������������������       �      ȼ"       ������J@�t�bh�hhK ��h��R�(KK�KK��h �Bh  ��k(/d@-����/c@������c@������a@��`@;��8�cP@2����"Z@j��F:lY@��-��-5@�5��X@������S@vb'vb'"@�k(���U@��h
�G@H�4H�4@��Gp_R@��h
�G@H�4H�4@��#���?���-��@                0����/@        ��#���?��/����?        ��#���?                        ��/����?        �YLg1R@'jW�v%D@H�4H�4@�P^CyO@%jW�v%D@H�4H�4@z�5��@�cp>'@        z�5��@0����/@        z�5��@��/����?                ��/����?        z�5��@                        �cp>@                ���-��@            �M@��|��<@H�4H�4@<��,��D@�cp>@        =��,��D@�cp>@        ��#�� @�cp>@        ��#�� @                        �cp>@        ��#��@@                Jp�}>@                z�5��@                        �cp>@        ��,���1@�cp>7@H�4H�4@|�5��(@�cp>7@H�4H�4@��#��@:l��F:2@H�4H�4@��#��@��/���@0#0# @��#��@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ��#�� @                        �cp>@0#0# @        �cp>@0#0#�?                0#0#�?        �cp>@                        0#0#�?        ��|��,@0#0#�?        ��On�(@                ��/����?0#0#�?                0#0#�?        ��/����?        ��#�� @0����/@        z�5��@                ��#�� @0����/@                ��/���@        ��#�� @��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                ;��,��@                ��#���?                ��#��@                <��,��$@                ��b:��*@                z�5��(@�]�ڕ�?@H�4H�4@�k(��"@�]�ڕ�?@0#0#@z�5��@�cp>�9@        z�5��@0����/#@        ��#���?0����/#@                ��/���@        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                        On��O0@                E�JԮD!@                ��/���@        z�5��@�cp>@0#0#@��#�� @�cp>@        ��#�� @                        �cp>@                �cp>@                �cp>@        ��#��@        0#0#@��#��@                                0#0#@z�5��@        0#0# @z�5��@                                0#0# @;��,��@�cp>7@H�4H�4(@z�5��@��/���.@        ��#�� @��/���.@        ��#���?��/���.@        ��#���?��/����?                ��/����?        ��#���?                        ���-��*@        ��#���?                ��#���?                ��#�� @��/���@H�4H�4(@        ���-��@H�4H�4@        �cp>@0#0#�?        �cp>@0#0#�?        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@                ��/����?0#0# @                0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?        ��#�� @��/����?vb'vb'"@��#���?        vb'vb'"@                H�4H�4@��#���?        H�4H�4@                0#0# @��#���?        0#0#�?                0#0#�?��#���?                ��#���?��/����?                ��/����?        ��#���?                d:��,&C@���-��:@#0#0F@��#��@@%jW�v%4@%S2%S27@�P^Cy?@��|��,@%S2%S27@�P^Cy?@���-��*@��8��8*@+�����;@鰑%@        |�5��8@��/���@        \Lg1��6@�cp>@        \Lg1��6@��/����?        �k(��2@��/����?        <��,��$@��/����?        ��#���?��/����?        ��#���?                        ��/����?        �k(��"@                ��#�� @                ��#��@��/����?        ��#��@                        ��/����?                ��/����?        ��#�� @��/����?                ��/����?        ��#�� @                z�5��@���-��@                ���-��@                ��/����?                �cp>@        z�5��@                z�5��@�cp>@��8��8*@��#�� @�cp>@��8��8*@        �cp>@        ��#�� @        ��8��8*@                �C=�C=@��#�� @        H�4H�4@��#�� @        0#0#�?��#�� @                                0#0#�?                ��+��+@��#���?                        ��/����?��+��+$@        ��/����?                        ��+��+$@��#�� @�cp>@        ��#�� @��/����?        ��#�� @��/����?        ��#�� @                        ��/����?                ��/����?                ��/���@        ;��,��@���-��@��-��-5@;��,��@��/����?        ;��,��@��/����?        ��#���?                ��#��@��/����?        ��#���?��/����?                ��/����?        ��#���?                z�5��@                        ��/����?                0����/@��-��-5@        0����/@��+��+@        0����/@0#0#�?        �cp>@                ��/����?0#0#�?        ��/����?                        0#0#�?                0#0#@                0#0#0@�k(��2@��On�8@ �q��V@�k(��2@��On�8@��)��)C@�k(��2@��On�8@��-��-5@��b:��*@��/����?��+��+@[Lg1��&@��/����?0#0#�?��#���?        0#0#�?��#���?                                0#0#�?;��,��$@��/����?                ��/����?        ;��,��$@                ��#�� @        0#0#@                0#0#@��#�� @                ;��,��@�e�_��7@0#0#0@��#���?��/���.@0#0#@        �cp>@0#0#@        ��/����?                ��/����?0#0#@                0#0#@        ��/����?        ��#���?��On�(@        ��#���?��/���@        ��#���?��/����?        ��#���?                        ��/����?                �cp>@                ��/����?                ��/����?                E�JԮD!@        ��#��@D�JԮD!@H�4H�4(@                ��+��+@��#��@D�JԮD!@�C=�C=@        E�JԮD!@��+��+@        ��/����?��+��+@                0#0#@        ��/����?0#0#�?                0#0#�?        ��/����?                ���-��@        ��#��@        0#0# @��#���?        0#0# @��#���?                                0#0# @z�5��@                                S2%S2%1@                H�4H�4@                �C=�C=,@                ������J@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��(hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKӅ�h��B(.         �                 ��V�?����R�?"      T���x}@       ;                 0%�z?�@r�L��?�       ��6@>q@       6                 �jE?>�����?R       Q(�\Sg`@       #                 ~`�� �r�~��?I       ���<T�]@       
                   ��?���/��?       �ټ�|�I@                        ���`?e��}�?       ��Se+@������������������������       �      ȼ       /����/#@       	                 P.�?֔fm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@                        p6��?Zg׬��?       B��o�,C@                           �?�)z� ��?       �\�<@                        `f��>�Q0TuJ�?       Ƀ�Я[5@                        @.��>f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?                        �ny?�����?
       L��o�g2@                        (��a?T�s�	�?       d���*@������������������������       �      ��       ���>��@                        @*��?�����?       �O��@������������������������       �               ��/����?������������������������       �      �<       ;��,��@                         P�J�?֗Z�	7�?       j~���@������������������������       �               z�5��@������������������������       �      �<       ��/����?                        �<��>      �<       ���-��@������������������������       �               ��/����?������������������������       �               0����/@                           \��?�FO���?       �ߌ$@                         �JV�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?!       "                 hf�?      �<       ��#�� @������������������������       �               z�5��@������������������������       �               ;��,��@$       %                 0��?l�E�B��?+       �]�ڕ�P@������������������������       �               ��/����?&       5                   ��?xҁ
_�?*       ����/�P@'       4                 �x? ?6��,�?       us���D@(       -                 �m۶?X���m>�?       0w��e�B@)       *                  �9��?��F¯?       �:.�=@������������������������       �        	       ;��,��4@+       ,                   E(�?h�j���?       ���z"@������������������������       �               ��/����?������������������������       �               ��#�� @.       /                 �b?B9�)\e�?       _���b @������������������������       �               ��/����?0       1                 �a{?�����?       �O��@������������������������       �               z�5��@2       3                 аZ(?bn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ȼ       ��/���@������������������������       �               |�5��8@7       8                 ��?��fm���?	       �0��z'@������������������������       �      ȼ       �cp>@9       :                 @� %?���/��?       @z$S��@������������������������       �               z�5��@������������������������       �               �cp>@<       m                 `8��?��S�4��?W       @�#)�a@=       Z                 ����?#S����?7       '���mU@>       M                 �Fq?x�ut��?%       ��R�I@?       L                 ��|�?�	>�S�?       ���FV%?@@       E                 P��?z1���?       �8���<@A       D                 8*��?)���?       y��uk1@B       C                 �:=�?��i�@M�?       ���wzb0@������������������������       �               ��/���.@������������������������       �      �<       ��#���?������������������������       �      �<       ��#���?F       K                 ��Z�?������?       ,�ǟf%@G       J                 pL��?�w��d��?       �0���s@H       I                 @Ͳ�?putee�?       Q9��@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?������������������������       �      м       ��/����?������������������������       �      ��       ��/���@������������������������       �               H�4H�4@N       W                  `s�?�x�I��?       ��]\3@O       V                 @$�?"3�Ҽ��?
       ����@,@P       Q                  ~��?&���
�?	       䡍�C&@������������������������       �               z�5��@R       S                 P�L�?����]L�?       N66�ͯ@������������������������       �               �cp>@T       U                 lh#s?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �      �<       �cp>@X       Y                 �J�?�o���?       o�9�F@������������������������       �               0#0#@������������������������       �               ��#���?[       \                 �-�?�fL�z��?       2r�%�A@������������������������       �               ��/����?]       j                 �jE?ܕ��+�?       <���@@^       c                 `���?��^��\�?       F��⋣=@_       b                 �؉�?�hK)�?
       �h��K�2@`       a                �3G�y?�����?       �O��@������������������������       �               ��/����?������������������������       �               ;��,��@������������������������       �               z�5��(@d       i                    �?4k�"O��?       �?<��*&@e       h                 �3�?j��H��?       v�I�@f       g                 p%�?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@������������������������       �               �cp>@������������������������       �               ��#��@k       l                 @�ԏ?v�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @n       }                  �ni?iV-���?        ԮiJ�`L@o       |                  1��?�ޱ��?       ��}��nD@p       s                 �;�?�_�t�#�?       �`�`Zy:@q       r                 �-�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@t       w                 0��?j��M�?       7B��	�2@u       v                 ��'�?      �<       �cp>'@������������������������       �               �cp>@������������������������       �               E�JԮD!@x       {                 �HQ�?���q���?       �:-ߩ�@y       z                  �ƫ?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �               z�5��@������������������������       �      ��       ��|��,@~       �                 ��=~?��h����?       ��[�/@       �                 @x��?�v�;B��?       ՟���	 @������������������������       �               H�4H�4@�       �                 ���?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 �TI�?|�G���?       ��%�|@������������������������       �               �cp>@�       �                  ��^�?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?�       �                 �WZ�?���Lq�?y       .e���h@�       �                 '�\?�~{U��?X       ��2�a@�       �                   �g�?��+�n��?4       a��]�U@������������������������       �               鰑%@�       �                 �I��?vAv����?/       @�J���R@�       �                 �U��>"����a�?       8It��B@�       �                 0�3�?������?       8u$Tml:@�       �                  ��?<9�)\e�?       _���b @������������������������       �               ;��,��@������������������������       �               �cp>@�       �                 е?H����?       �����^2@������������������������       �               H�4H�4@�       �                 �Tʡ?^�Ua4�?
       >
�#W�.@�       �                 p��?�i^�c�?       �D9�V$@�       �                  _�?�@����?       ���a�@������������������������       �               ��/����?������������������������       �               0#0#@������������������������       �      �<       ;��,��@������������������������       �      ��       ;��,��@�       �                    �?���3�?       ���(+�%@�       �                 P�T�?���/��?       U��7�@������������������������       �               ��/����?�       �                  �/�?\n����?       � ��w<@������������������������       �               z�5��@�       �                 �vA�?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      Լ       �cp>@�       �                 `7h�?�f���\�?       h�Lv6.C@�       �                      W�йT�?       �|Pp�L=@�       �                 0��?�4�fP�?	       V���-@�       �                    �?0��~d��?       7E���*@�       �                  pjS�?���mf�?       毠�?b@������������������������       �      �<       ��/���@������������������������       �               0#0#�?������������������������       �               D�JԮD!@������������������������       �      �<       ��#���?�       �                 P� �?���d��?	       ��GQ�-@�       �                 @E��?�@G���?       hu��@������������������������       �               0����/@�       �                 h�R?z��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?�       �                 pj��?X�ih�<�?       ��
@������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?�       �                  `��?H��aB��?       ����"@�       �                 �Ծ�?      �<       ;��,��@������������������������       �               ��#���?������������������������       �               ��#��@�       �                  `s�?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@�       �                    �?�{�JѠ?$       P���L@�       �                 ��
�?      �<       �ڬ�ڬD@������������������������       �               H�4H�4@������������������������       �               ��)��)C@�       �                 ��>�?�q����?
       Qz�i0@�       �                 ���?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 p'v�?      �<       ��8��8*@������������������������       �               0#0#�?������������������������       �               H�4H�4(@�       �                   �0�?Ԥ��Q��?!       �X0�K@�       �                 @��?�E���?       �|����4@�       �                 pdJ�?�� ��?       rp� k@������������������������       �               0#0# @������������������������       �      �<       ��/���@�       �                 �!�?��(v��?	       �A�s(.@������������������������       �               ��+��+$@�       �                 Į�?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?������������������������       �               B�A�@@�t�bh�hhK ��h��R�(KK�KK��h �B�  g:��,&c@�����d@�؉��Ic@Jy�5�_@��|��\@=�C=�C?@�GpAV@鰑E@        ����bzU@�-����@@        ��b:��:@��On�8@        ��#���?��On�(@                /����/#@        ��#���?�cp>@        ��#���?                        �cp>@        
�#���9@��On�(@        ��#��0@�cp>'@        ��#��0@0����/@        ��#���?��/����?        ��#���?                        ��/����?        �P^Cy/@�cp>@        z�5��(@��/����?        ���>��@                ;��,��@��/����?                ��/����?        ;��,��@                z�5��@��/����?        z�5��@                        ��/����?                ���-��@                ��/����?                0����/@        �k(��"@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                z�5��@                ;��,��@                    �M@D�JԮD!@                ��/����?            �M@��/���@        Ey�5A@��/���@        Dy�5A@��/���@        ���>��<@��/����?        ;��,��4@                ��#�� @��/����?                ��/����?        ��#�� @                ;��,��@�cp>@                ��/����?        ;��,��@��/����?        z�5��@                ��#�� @��/����?                ��/����?        ��#�� @                        ��/���@        |�5��8@                z�5��@D�JԮD!@                �cp>@        z�5��@�cp>@        z�5��@                        �cp>@        e:��,&C@;l��F:R@=�C=�C?@��,���A@�+Q��B@��8��8*@<��,��$@��|��<@#0#0&@��#�� @�cp>7@H�4H�4@��#�� @�cp>7@H�4H�4@��#�� @��/���.@        ��#���?��/���.@                ��/���.@        ��#���?                ��#���?                        ��/���@H�4H�4@        ��/���@H�4H�4@        ��/����?H�4H�4@                H�4H�4@        ��/����?                ��/����?                ��/���@                        H�4H�4@��#�� @�cp>@��+��+@���>��@�cp>@0#0#�?���>��@�cp>@0#0#�?z�5��@                ��#���?�cp>@0#0#�?        �cp>@        ��#���?        0#0#�?                0#0#�?��#���?                        �cp>@        ��#���?        0#0#@                0#0#@��#���?                {�5��8@D�JԮD!@0#0# @        ��/����?        z�5��8@���-��@0#0# @z�5��8@0����/@        ��,���1@��/����?        ;��,��@��/����?                ��/����?        ;��,��@                z�5��(@                ���>��@��/���@        z�5��@��/���@        z�5��@��/����?                ��/����?        z�5��@                        �cp>@        ��#��@                        ��/����?0#0# @        ��/����?                        0#0# @z�5��@����z�A@vb'vb'2@z�5��@��/���>@�C=�C=@z�5��@Nn��O0@�C=�C=@        ��/����?H�4H�4@        ��/����?                        H�4H�4@z�5��@��|��,@0#0#�?        �cp>'@                �cp>@                E�JԮD!@        z�5��@�cp>@0#0#�?        �cp>@0#0#�?                0#0#�?        �cp>@        z�5��@                        ��|��,@                0����/@#0#0&@        ��/����?�C=�C=@                H�4H�4@        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/���@0#0#@        �cp>@                ��/����?0#0#@                0#0#@        ��/����?        
�#���9@z%jW�vH@/��+��^@�#���9@h
��F@���~�gR@
�#���9@��]�ڕE@S2%S2%1@        鰑%@        
�#���9@Pn��O@@S2%S2%1@������3@鰑%@�C=�C=@�P^Cy/@��/���@�C=�C=@;��,��@�cp>@        ;��,��@                        �cp>@        ;��,��$@��/����?�C=�C=@                H�4H�4@;��,��$@��/����?0#0#@;��,��@��/����?0#0#@        ��/����?0#0#@        ��/����?                        0#0#@;��,��@                ;��,��@                ��#��@���-��@        ��#��@��/���@                ��/����?        ��#��@��/����?        z�5��@                ��#���?��/����?        ��#���?                        ��/����?                �cp>@        z�5��@h
��6@��+��+$@��#���?0����/3@vb'vb'"@��#���?��On�(@0#0#�?        ��On�(@0#0#�?        ��/���@0#0#�?        ��/���@                        0#0#�?        D�JԮD!@        ��#���?                        ���-��@0#0# @        �cp>@0#0# @        0����/@                ��/����?0#0# @                0#0# @        ��/����?                ��/����?H�4H�4@                H�4H�4@        ��/����?        ;��,��@�cp>@0#0#�?;��,��@                ��#���?                ��#��@                        �cp>@0#0#�?                0#0#�?        �cp>@                ��/����?�C=�C=L@                �ڬ�ڬD@                H�4H�4@                ��)��)C@        ��/����?�A�A.@        ��/����?0#0# @        ��/����?                        0#0# @                ��8��8*@                0#0#�?                H�4H�4(@        0����/@Z��Y��H@        0����/@0#0#0@        ��/���@0#0# @                0#0# @        ��/���@                ��/����?�C=�C=,@                ��+��+$@        ��/����?0#0#@                0#0#@        ��/����?                        B�A�@@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ���~hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKᅔh��B81         p                 pS�?\�uɪ4�?)      ���~}@       e                 ��c�?��#��?�       �^[" p@       d                 �+��?G�Nܚd�?�       ���o��m@                        0��Q?�������?�       d
^Q�
m@                        � �l?�O-r��?       �.w��e9@                         @�a�?�^�#΀�?       O�{��A5@       
                 P�_?��٤ݸ?       ��<5�84@       	                 0��>f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �        	       D�JԮD1@������������������������       �      �<       ��#���?������������������������       �               ��#��@       7                 P �s?�ګ!uJ�?~       �$O���i@       4                 ���?H�sBB�?E       ��C�o]@       )                  p�:?675��5�?C       ��o<u\@       &                 p���?0eI�LX�?3       :�~��W@                        )DW?x%����?1       n�ZDV@                        �U���������?$       8nҟ��O@                          �P�?�����?
       �O��8@                        �7�<?�hK)�?       �h��K�2@                        �Π+?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �      ��       ��b:��*@                        �e�O?���/��?       @z$S��@������������������������       �               �cp>@������������������������       �               z�5��@������������������������       �      ��       ������C@       %                 �(+�?\]���?       ��29@       $                 �=y?���/��?
       �[[�.�1@        !                 � ��?4=�%�?	       t=�x�-@������������������������       �               ��/���@"       #                 p��h?�PJo�x�?       U|qt�&@������������������������       �               z�5��@������������������������       �               0����/@������������������������       �      ȼ       z�5��@������������������������       �      ��       ���>��@'       (                 �L+�?E#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @*       +                 ��,b?r��3�?       ���(+�5@������������������������       �               ��#��@,       1                    �?rQ��?       �s�=�1@-       .                 0�?���3�?	       ���(+�%@������������������������       �               ��/���@/       0                 �iDe?�)z� ��?       ~�\�@������������������������       �               ��#��@������������������������       �      ȼ       �cp>@2       3                  �P��?      �<       ���-��@������������������������       �               ��/����?������������������������       �               0����/@5       6                �OORp?��fm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@8       U                 0�`�?7�C8J�?9       ��nDLV@9       F                 ����?@�\�4b�?#       _���IG@:       ;                 ��?B�,��y�?       ��V6@������������������������       �               ��/����?<       C                 �K��?��7m�?       �(�+4@=       >                  ;��?�HU����?       !��N��%@������������������������       �               z�5��@?       @                 �nF�?ʔfm���?       ��Z�N@������������������������       �               0����/@A       B                ��W�y?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @D       E                 ����?��j���?       ���z"@������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?G       H                  �\�?�_�ѡ��?       �`��|8@������������������������       �               �cp>@I       P                  �!�?p1Y�RM�?       g�h4�2@J       O                 ��(�?�n�l���?       ���5F'@K       N                 `s5�?�}	;	�?       vK�>4%@L       M                 ��Z�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               ��/���@������������������������       �      �<       ��#���?Q       T                 ��=�?�_�A�?       肵�e`@R       S                 ����?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               z�5��@V       [                  Ϳ�?^<��;�?       �z�W�NE@W       X                 �Gn�?~�����?       �4^$4�#@������������������������       �               �cp>@Y       Z                 �5W�?�����?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?\       c                    �?��b���?       ��N�e@@]       `                  @?��?j-�=H�?       "<��R,@^       _                 8��H?,Lj����?       ���T�@������������������������       �               z�5��@������������������������       �               0#0#�?a       b                 ��<�?h��H��?       v�I�@������������������������       �               ��/���@������������������������       �      ��       z�5��@������������������������       �      ��       �k(��2@������������������������       �     ��       �C=�C=@f       i                 ����?B!A_!�?       E����0@g       h                  Џ~�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@j       k                  ���?�L����?       Yk���>)@������������������������       �               ��#���?l       m                  I�4?�F���?       :�.�-'@������������������������       �      ��       E�JԮD!@n       o                 ����?j%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?q       �                 �{��?x����Z�?�       "�`a�j@r       y                 ��Ǆ?��N:��?8       >&�L�V@s       x                 e�h?���_�?       ���e��#@t       w                 ��~?��b�}�?       ���\�@u       v                 �ǽv?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �               0����/@z       �                 ��Ҧ?�v���E�?0       ��=XxT@{       |                   �?,��,��?       ����J@������������������������       �               �C=�C=<@}       �                  �׽�?�۞�ڳ�?       ;����9@~                         ���?֞�z�F�?       �]!_��5@������������������������       �               ��/����?�       �                 (a�?�Y�����?       ���o]5@�       �                    �?xT �+��?       ��>Y��@�       �                  �Ԧ�?Δfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               0#0# @�       �                  �6��?��(v��?
       �A�s(.@������������������������       �               #0#0&@�       �                 �j%?����|e�?       �z �B�@������������������������       �               0#0# @�       �                 �.�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ȼ       z�5��@�       �                 ��
�?�
͎�y�?       ��ڦ��:@�       �                 P㕸?���`�?       ��
�Me@������������������������       �               ��/���@�       �                 ���?�3`���?       .�r��@������������������������       �               ��#���?�       �                 ���?���`p��?       �����@������������������������       �               0#0#�?�       �                 �b'�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 �$I�??�	,�?       >0�1b3@������������������������       �               ��8��8*@�       �                 xr��?z��`p��?       �����@������������������������       �               0#0# @�       �                 �ޥg?|�G���?       ��%�|@������������������������       �               0#0#�?�       �                 �z��?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?�       �                 ����?xr2:���?U       ǽ�v_@�       �                 ���?��E���?K       �e?C6�[@�       �                    �?��.���?       ܪU=>@�       �                   ��?x���ߡ�?
       г"�-@������������������������       �               ��/���@�       �                 (�0m?�ݛ��4�?       #�V�%�%@�       �                 �*��?A��X�&�?       �6��	�@�       �                 �?Pw?& k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      �<       ��/���@�       �                 �`	�?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?������������������������       �               H�4H�4@�       �                 0�y?�Tu��?       ����.@������������������������       �               ��#���?������������������������       �      ��       ��|��,@�       �                 �Է�?�h_���?9       ົ��_T@�       �                 �Y�?(g���?       ��+���*@�       �                 `�;�?�FO���?
       �ߌ$@�       �                  �я�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @�       �                     �?      �<       ���>��@������������������������       �               ��#���?������������������������       �               z�5��@������������������������       �               H�4H�4@�       �                  V��?��Fy��?-       �=��Q@�       �                  �fq?��K=^�?'       ����N@�       �                  �d%�?\�0a��?       ���*X�A@�       �                  �6��?�{��?       ����*>@�       �                 `��?���i�?       7����s7@�       �                 �I��?�C1���?       "@��9l4@�       �                 h��1?l��H��?       v�I�@�       �                ��?��?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@������������������������       �               �cp>@�       �                  ��??L��~d��?       7E���*@�       �                 �9/�?�֪u�_�?       ��?�8@������������������������       �               ��/���@�       �                 _%?z�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       ��/���@�       �                 i��?ln����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               ���-��@�       �                  �{��?jutee�?       Q9��@������������������������       �               0#0#�?�       �                 �p�?|�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 7��?���@��?       �<��9@������������������������       �               #0#06@������������������������       �      �<       �cp>@�       �                  ��d�?w�;B��?       ՟���	 @�       �                  �g<�?|��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               ��+��+@�       �                 0���?      �<
       �C=�C=,@������������������������       �               0#0#�?������������������������       �        	       ��8��8*@�t�bh�hhK ��h��R�(KK�KK��h �B  ����bze@[�ڕ��d@D�A�`@�5��P>b@�e�_��W@�C=�C=,@�}��a@鰑U@#0#0&@�}��a@鰑U@0#0#@z�5��@/����/3@        ��#�� @/����/3@        ��#���?0����/3@        ��#���?��/����?                ��/����?        ��#���?                        D�JԮD1@        ��#���?                ��#��@                YUUUU5a@Qn��OP@0#0#@�k(���U@��|��<@0#0# @����bzU@�cp>�9@0#0# @���khS@��On�(@0#0# @f:��,&S@��On�(@        Np�}N@��/���@        ;��,��4@��/���@        ��,���1@��/����?        ��#��@��/����?        ��#��@                        ��/����?        ��b:��*@                z�5��@�cp>@                �cp>@        z�5��@                ������C@                ��#��0@E�JԮD!@        �k(��"@D�JԮD!@        z�5��@E�JԮD!@                ��/���@        z�5��@0����/@        z�5��@                        0����/@        z�5��@                ���>��@                ��#���?        0#0# @��#���?                                0#0# @��#�� @���-��*@        ��#��@                ��#��@���-��*@        ��#��@���-��@                ��/���@        ��#��@�cp>@        ��#��@                        �cp>@                ���-��@                ��/����?                0����/@        ��#���?�cp>@        ��#���?                        �cp>@        �}�\I@;l��F:B@0#0# @������3@�cp>�9@0#0#�?��b:��*@D�JԮD!@                ��/����?        ��b:��*@���-��@        ;��,��@�cp>@        z�5��@                ��#�� @�cp>@                0����/@        ��#�� @��/����?                ��/����?        ��#�� @                ��#�� @��/����?        ��#�� @                        ��/����?        z�5��@D�JԮD1@0#0#�?        �cp>@        z�5��@�cp>'@0#0#�?��#���?/����/#@0#0#�?        0����/#@0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                ��/���@        ��#���?                ;��,��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        z�5��@                �P^Cy?@鰑%@0#0#�?z�5��@���-��@                �cp>@        z�5��@��/����?        z�5��@                        ��/����?        )�����;@��/���@0#0#�?�k(��"@��/���@0#0#�?z�5��@        0#0#�?z�5��@                                0#0#�?z�5��@��/���@                ��/���@        z�5��@                �k(��2@                                �C=�C=@��#�� @�cp>'@H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@��#�� @鰑%@        ��#���?                ��#���?鰑%@                E�JԮD!@        ��#���?��/����?                ��/����?        ��#���?                �#���9@����z�Q@����]@���>��@:l��F:2@2#0#P@��#�� @���-��@0#0#�?��#�� @��/����?0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?        ��#�� @                        0����/@        ;��,��@�cp>'@O��N��O@��#��@0����/@#0#0F@                �C=�C=<@��#��@0����/@0#0#0@��#���?0����/@0#0#0@        ��/����?        ��#���?��/���@0#0#0@��#���?�cp>@0#0# @��#���?�cp>@        ��#���?                        �cp>@                        0#0# @        ��/����?�C=�C=,@                #0#0&@        ��/����?H�4H�4@                0#0# @        ��/����?0#0#�?        ��/����?                        0#0#�?z�5��@                ��#���?���-��@��)��)3@��#���?0����/@0#0# @        ��/���@        ��#���?��/����?0#0# @��#���?                        ��/����?0#0# @                0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                ��/����?S2%S2%1@                ��8��8*@        ��/����?0#0#@                0#0# @        ��/����?0#0# @                0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?�k(��2@b#6�aJ@�;�;K@�k(��2@c#6�aJ@��+��+D@��#��@h
��6@0#0#@z�5��@��/���@0#0#@        ��/���@        z�5��@��/���@0#0#@z�5��@��/���@0#0#�?��#���?��/���@        ��#���?                        ��/���@        ��#�� @        0#0#�?��#�� @                                0#0#�?                H�4H�4@��#���?��|��,@        ��#���?                        ��|��,@        ���>��,@��/���>@wb'vb'B@�k(��"@��/����?H�4H�4@�k(��"@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ���>��@                ��#���?                z�5��@                                H�4H�4@;��,��@�_��e�=@B�A�@@;��,��@��|��<@��8��8:@;��,��@�cp>�9@0#0#@;��,��@�e�_��7@0#0#�?;��,��@D�JԮD1@0#0#�?z�5��@On��O0@0#0#�?z�5��@��/���@        z�5��@��/����?                ��/����?        z�5��@                        �cp>@                ��On�(@0#0#�?        0����/@0#0#�?        ��/���@                ��/����?0#0#�?        ��/����?                        0#0#�?        ��/���@        ��#�� @��/����?        ��#�� @                        ��/����?                ���-��@                ��/����?H�4H�4@                0#0#�?        ��/����?0#0# @        ��/����?                        0#0# @        �cp>@#0#06@                #0#06@        �cp>@                ��/����?�C=�C=@        ��/����?0#0# @                0#0# @        ��/����?                        ��+��+@                �C=�C=,@                0#0#�?                ��8��8*@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJCLUhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKׅ�h��B/         v                  �?�I�)�T�?'      1l�?ɂ}@       a                 �T�x?��� ��?�       z�S:�p@       4                 p��v?Z_�h��?t       ZG䁭h@       -                  |v?>��m"�?A       MH�3f�Y@       (                 �jE?v:R����?9       ~bݻ��V@                        �U���̍��b�?1       T�f\T@                        ���?��U>��?       �Y�^�3@                           �?&r��lB�?       ��%��t/@	                        0��j?Bǵ3���?       �q�ͨ�@
                          B�?r@ȱ��?       nm���S@������������������������       �      ��       0����/@������������������������       �               ��#���?������������������������       �               ��#�� @                        �Q�?Ȕfm���?       ��Z�N@������������������������       �               0����/@                        h�-V?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @                         �g<�?      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@       '                 ܙ?������?!       @{;���N@                         y��?��(���?       �ټ�|=@                        �QZ?X ����?       2
C>�5@������������������������       �               ��#��0@                        �>�#?�d�$���?       �T�f@������������������������       �               z�5��@                        VV?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?       &                    �?̔fm���?       ��Z�N@        !                 �_�?d%@�"�?       ��[�@������������������������       �               �cp>@"       #                 bq(?Zn����?       � ��w<@������������������������       �               ��#���?$       %                 Њ�8?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��/����?������������������������       �               ���b:@@)       ,                 ����?Q��?       �s�=�!@*       +                  �{��?h�r{��?       e�6� @������������������������       �               ���-��@������������������������       �               ��#���?������������������������       �               ��#���?.       /                 pA}?��O-r��?       �.w��e)@������������������������       �               �cp>@0       3                 �I?h��H��?       v�I�@1       2                 (`��?d%@�"�?       ��[�@������������������������       �      �<       ��/���@������������������������       �               ��#�� @������������������������       �               ��#���?5       ^                 4��?沂?�n�?3       l�����W@6       M                 P�>�?@�����?1       ?�h�\V@7       8                   ��?8����?"       *�լ�^N@������������������������       �               ��/���.@9       J                 ����?Dv�P�g�?       z�	2�F@:       I                  �]?d9��;3�?       �ll�D@;       <                 �5W�?��9��8�?       �+M��C@������������������������       �               ;��,��@=       D                  �Q�?`ҭ�?��?       b��� A@>       A                  �\�?e��}�?       ��Se;@?       @                 �8�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?B       C                 �L0?���gN�?       �F���9@������������������������       �               ��#���?������������������������       �               �e�_��7@E       F                 �Dָ?���q���?       �:-ߩ�@������������������������       �               �cp>@G       H                    �?�zœ���?       IG���t@������������������������       �               0#0#�?������������������������       �               z�5��@������������������������       �               ��#���?K       L                  ����?      �<       ;��,��@������������������������       �               ��#��@������������������������       �               ��#���?N       W                    �?�\�����?       ���I�<@O       V                 �j%?fQ ����?
       +�_ݗ�3@P       S                 0�!�?����>��?       �>@a@.@Q       R                 ���?�"6Aq�?       )$�B"@������������������������       �               ��#�� @������������������������       �               �C=�C=@T       U                 0I��?x�G���?       '5L�`�@������������������������       �               �cp>@������������������������       �               H�4H�4@������������������������       �               0����/@X       ]                 h��1?�Ϟi�?       ��ؠ�!@Y       Z                 @�#�?Ny��]0�?       ���y"@������������������������       �               0#0#@[       \                  ���?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               �cp>@_       `                 ����?      �<       ��+��+@������������������������       �               0#0# @������������������������       �               H�4H�4@b       k                    �?Z�����?)       3�E���P@c       j                 Ț_c?<�y;��?       �\�K�?@d       e                  ��^�?�=�Sο?       ����<@������������������������       �               ������3@f       g                 _%?L���'0�?       �C�� T"@������������������������       �               ;��,��@h       i                 ���?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               H�4H�4@l       o                 ȏ�B?��!�j�?       ��}K%�A@m       n                 @�?      �<       �k(���5@������������������������       �        	       ��#��0@������������������������       �               ;��,��@p       q                 �5�?0�Z�K��?	       X��Q�+@������������������������       �               ��+��+@r       s                 �oW�?�����?       �v�qp�!@������������������������       �               H�4H�4@t       u                  0B�?�֪u�_�?       ��?�8@������������������������       �               0����/@������������������������       �               0#0#�?w       �                 �6Sz?��� ;-�?�       �����i@x       �                   s��?���2���?\       ���]xa@y       �                 �se?��,��?!       #�Gn�J@z       �                 ���@?ĸ�qA��?       �����5@{       �                 ����?$Й����?       �3�N0@|       �                  �g<�?d����?	       P	K��,@}       �                 ����?`�s�	�?       d���*@~       �                 P6��?\����?       P	K��@       �                 Ш��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ��       ;��,��@������������������������       �      ȼ       z�5��@������������������������       �      ȼ       ��/����?�       �                 d[�?v�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                    �?      �<       0����/@������������������������       �               ��/����?������������������������       �               �cp>@�       �                 �&^�?�DW��?       �˅k
@@�       �                 ��:�?�Tu��?       ����.@������������������������       �      ȼ       �cp>'@�       �                 PW�?Ȕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?�       �                 �
�k?�P�`B�?       �F�N@�0@�       �                 PFe�?��[����?	       Hl�_A+@�       �                 @?�����?       �v�qp�!@�       �                 �$I�?�@����?       ���a�@������������������������       �               ��/����?������������������������       �               0#0#@������������������������       �      ��       ��/���@������������������������       �      ȼ       0����/@������������������������       �               H�4H�4@�       �                 P�/|?
��U�?;       �LN�U@�       �                 ����?���f��?       ��>�BzE@�       �                  �~��?Py��]0�?       ���y"8@������������������������       �               ��/����?�       �                 ��?��q��?       �?8��7@������������������������       �               �C=�C=@�       �                 0�rM?f�q����?       O�Q*s�/@�       �                   ��?�n���k�?	       3��&�*@������������������������       �               H�4H�4@�       �                  ���?X�ih�<�?       ��
@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                 0\?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?�       �                    �?T����?       �|�c�2@�       �                 �U�,?�3`���?       .�r�� @������������������������       �               H�4H�4@�       �                  �5�?��b�}�?       ���\�@������������������������       �               ��#�� @�       �                  �{��?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?�       �                 �"�?^H-����?       p�c#��%@�       �                   �0�?& k�Lj�?       �q��l}@������������������������       �               ��/����?�       �                  0Y��?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ��       H�4H�4@�       �                 `���?R����?       {�Y���E@������������������������       �               0����/@�       �                  /U�?�w̙��?       ����iC@������������������������       �               ��/����?�       �                 �D���ݹ�7�?       e��1tB@�       �                 p��?z�����?       �4^$4�#@�       �                 K��?��Z�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@������������������������       �               0����/@�       �                 �\��?xļm�6�?       ԯ�I;@�       �                 �lw?�&t�ׁ�?       3�1!�4@�       �                 ���?�#Vn\��?       H�~B�2@������������������������       �      ��       �A�A.@�       �                 ���?���`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      ȼ       ��/����?�       �                 ��H�?��G9�?       ���=A@�       �                    �?r�T���?       ��e[�&@�       �                 PU��?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               0#0#�?������������������������       �               H�4H�4@�       �                  �G�?�K���?.       zz=��P@�       �                   ���?      �<$       �˷|˷I@������������������������       �               0#0#�?������������������������       �        #       k�6k�6I@�       �                 `���?xq����?
       Qz�i0@������������������������       �               ��/����?������������������������       �      �<	       �A�A.@�t�b�T!     h�hhK ��h��R�(KK�KK��h �B(  �����c@鰑Nc@�6k�6�c@Gy�5a@>�cp�W@B�A�@@�#����U@h
��V@��-��-5@j1��tVQ@�-����@@        ��#��P@�e�_��7@        ���b:P@D�JԮD1@        �k(��"@鰑%@        ;��,��@鰑%@        z�5��@0����/@        ��#���?0����/@                0����/@        ��#���?                ��#�� @                ��#�� @�cp>@                0����/@        ��#�� @��/����?                ��/����?        ��#�� @                ��#��@                ��#���?                z�5��@                �>��nK@���-��@        \Lg1��6@���-��@        <��,��4@��/����?        ��#��0@                ��#��@��/����?        z�5��@                ��#���?��/����?                ��/����?        ��#���?                ��#�� @�cp>@        ��#�� @��/���@                �cp>@        ��#�� @��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                        ��/����?        ���b:@@                ��#�� @���-��@        ��#���?���-��@                ���-��@        ��#���?                ��#���?                z�5��@0����/#@                �cp>@        z�5��@��/���@        ��#�� @��/���@                ��/���@        ��#�� @                ��#���?                �k(��2@[�v%jWK@��-��-5@�k(��2@Z�v%jWK@0#0#0@��#��0@��]�ڕE@0#0#�?        ��/���.@        ��#��0@�a#6�;@0#0#�?ZLg1��&@�a#6�;@0#0#�?;��,��$@�a#6�;@0#0#�?;��,��@                ;��,��@�a#6�;@0#0#�?��#�� @��On�8@        ��#���?��/����?        ��#���?                        ��/����?        ��#���?�e�_��7@        ��#���?                        �e�_��7@        z�5��@�cp>@0#0#�?        �cp>@        z�5��@        0#0#�?                0#0#�?z�5��@                ��#���?                ;��,��@                ��#��@                ��#���?                ��#�� @�cp>'@�A�A.@��#�� @��/���@��+��+$@��#�� @�cp>@��+��+$@��#�� @        �C=�C=@��#�� @                                �C=�C=@        �cp>@H�4H�4@        �cp>@                        H�4H�4@        0����/@                ��/���@��+��+@        ��/����?��+��+@                0#0#@        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@                        ��+��+@                0#0# @                H�4H�4@4��tSH@���-��@H�4H�4(@��b:��:@��/����?H�4H�4@��b:��:@��/����?        ������3@                ���>��@��/����?        ;��,��@                ��#�� @��/����?        ��#�� @                        ��/����?                        H�4H�4@�k(���5@0����/@vb'vb'"@�k(���5@                ��#��0@                ;��,��@                        0����/@vb'vb'"@                ��+��+@        0����/@0#0#@                H�4H�4@        0����/@0#0#�?        0����/@                        0#0#�?�k(���5@�_��e�M@R`F`�_@�k(���5@F�)�BM@����M@��b:��*@�]�ڕ�?@0#0# @z�5��(@��/���@0#0#�?z�5��(@�cp>@0#0#�?z�5��(@��/����?        z�5��(@��/����?        z�5��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ;��,��@                z�5��@                        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?        0����/@                ��/����?                �cp>@        ��#���?�e�_��7@�C=�C=@��#���?��|��,@                �cp>'@        ��#���?�cp>@                �cp>@        ��#���?                        /����/#@�C=�C=@        0����/#@0#0#@        0����/@0#0#@        ��/����?0#0#@        ��/����?                        0#0#@        ��/���@                0����/@                        H�4H�4@��#�� @���-��:@~˷|˷I@z�5��@/����/#@�A�A>@        ��/���@��+��+4@        ��/����?                �cp>@��+��+4@                �C=�C=@        �cp>@��8��8*@        ��/����?H�4H�4(@                H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@        ��/����?0#0#�?        ��/����?                        0#0#�?z�5��@�cp>@��+��+$@��#�� @��/����?0#0#@                H�4H�4@��#�� @��/����?0#0#�?��#�� @                        ��/����?0#0#�?        ��/����?                        0#0#�?��#���?��/���@H�4H�4@��#���?��/���@                ��/����?        ��#���?��/����?        ��#���?                        ��/����?                        H�4H�4@;��,��@D�JԮD1@��-��-5@        0����/@        ;��,��@��On�(@��-��-5@        ��/����?        ;��,��@鰑%@��-��-5@z�5��@���-��@        z�5��@��/����?                ��/����?        z�5��@                        0����/@        ��#�� @��/���@��-��-5@        �cp>@S2%S2%1@        ��/����?S2%S2%1@                �A�A.@        ��/����?0#0# @        ��/����?                        0#0# @        ��/����?        ��#�� @��/����?0#0#@��#�� @��/����?0#0#�?��#�� @��/����?                ��/����?        ��#�� @                                0#0#�?                H�4H�4@        ��/����?D�A�P@                �˷|˷I@                0#0#�?                k�6k�6I@        ��/����?�A�A.@        ��/����?                        �A�A.@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ���hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK텔h��B�3         �                  ���?��	��M�?(      �bw�>t}@       Q                  �?���ɮ�?�       @���p@                         `���?K}����?^       �8�	zb@                         �x��?ʔfm���?       ��Z�N@������������������������       �               ��#�� @                        >^�l?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/���@	       8                 `%�7?_�Y@��?Y       �a�5	a@
                        P�`S?���-��?@       j�ޡ��X@                        ���U?h����?       ��x��A@                       h��\<?& k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      �<       ��/���@                         ����?�	�� ��?       A�x��>@������������������������       �               �#���9@                        �j?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?                         �_�?~���B��?(       	U��d�O@                        `s5�?��;�1�?
       �$�S՞1@������������������������       �               z�5��@                        �\͵?�4�fP�?       V���-@                        ����?�F���?       :�.�-'@                        �f�n?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               0����/#@                        @���?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?        +                 NK�X?���O�!�?       ���!��F@!       &                 PNs�?J��@���?       |�m�c1@"       #                  �ޖ?\����?       P	K��@������������������������       �               ��#��@$       %                 h��?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @'       (                 ����?����]L�?       N66�ͯ#@������������������������       �               �cp>@)       *                 PPp�?�J���?       ��*]Y@������������������������       �               ��#�� @������������������������       �               0#0# @,       /                 ���`?�Z�!���?       ��e`��<@-       .                 P&�s?
4=�%�?       �(J��@������������������������       �               ��#�� @������������������������       �               �cp>@0       5                 ��?��sx�?       �iۍѧ7@1       2                 py?�d�$���?       �T�f$@������������������������       �               ���>��@3       4                 �U��>`%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?6       7                 p'v�?      �<	       ��b:��*@������������������������       �               ��#���?������������������������       �               {�5��(@9       L                 0�2�?��˵��?       �KD��B@:       K                 �V:�?�Q&�Q�?       ������>@;       H                  ��d�?�u�N��?       ������=@<       E                  �_�?��'1��?       %�B��;@=       >                 @F��#�8b�?       �Ǣ�98@������������������������       �      ��
       D�JԮD1@?       @                 �\8?�`@s'��?       Ei_y,*@������������������������       �               �cp>@A       B                  ]P?Ȕfm���?       ��Z�N@������������������������       �               ��#���?C       D                 ��K?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?F       G                 �2OF?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@I       J                 � ��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               0#0#�?M       P                  �9��?l����1�?       ��;9�@N       O                 ���?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?������������������������       �               z�5��@R       �                 p��{?�#��|��?H       ��Y���^@S       �                 �c6�?��6x��?7       �)����W@T       u                 P7&E?�k�b��?1       ��U�K4T@U       j                 ��?H ��`��?       j�@��tH@V       _                 �&�?�~�1|�?       zi0���@@W       X                 �=�?����� �?       ��'���(@������������������������       �               0#0# @Y       \                 0u�?�FO���?       �ߌ$@Z       [                 ���?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?]       ^                 ���?      �<       ;��,��@������������������������       �               ��#�� @������������������������       �               z�5��@`       g                  ���?,Iz�9��?       ��[5@a       f                    �?�O
�*Q�?
       �͉V�M2@b       c                 @�C�?d�r{��?       e�6� @������������������������       �               0����/@d       e                 �U�,?b%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               鰑%@h       i                 ����?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?k       t                 0pS�?��v���?	       ��A蒇.@l       m                 p���?��q��?       ��4rz(@������������������������       �               H�4H�4@n       o                 �b'�?޺W�w��?       �'DQm"@������������������������       �               ;��,��@p       s                 @8��?u�T���?       ��e[�&@q       r                  P�"�?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �               H�4H�4@v       y                  "�?�,2��?       ���܎�?@w       x                  H(B�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@z                         �a�?�vQ�(�?       -�t�f�;@{       |                 ���?����x�?       
�ra6�:@������������������������       �               ��On�8@}       ~                 xQ}�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0#�?�       �                  X3�?�)w�q�?       ��|��-@�       �                 xs�?���mf�?       毠�?b@������������������������       �               0#0#�?������������������������       �      �<       ��/���@������������������������       �      ��       ��+��+$@�       �                 �p�?�)�n�?       �b�}{.;@������������������������       �      ��       #0#06@�       �                 �s�?�@����?       ���a�@�       �                 `���?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       H�4H�4@�       �                 p��{?�<c�+�?�       ԫn�?�i@�       �                 `{6�?�h��*�?]       1m��w|a@�       �                 ���@?AK��`^�?R       .� ���]@�       �                 �J�?�����?;       ǲ9�V@�       �                  ���?D�X���?/       Ҝ����Q@�       �                 `8X?��T[�?+       �dv�mP@�       �                 `s5�?��|��?       ���ĺw@������������������������       �               ��#�� @������������������������       �               0����/@�       �                   �0�?���w���?&       �c*�GlM@�       �                 @�C�?�����?
       �����1@�       �                 X��?�zœ���?       IG���t @������������������������       �               z�5��@������������������������       �               0#0# @������������������������       �               �k(��"@�       �                 @��>x����?       ��P ��D@������������������������       �               ��#��@�       �                    �?�ʍ+F_�?       `��B@�       �                 �a�?��h!��?       Z�v%jW;@�       �                 ��N�?��Ӭ%�?       ޅ��p3@�       �                  ���?�C=+��?
       b��T|0@�       �                 ��?L�j���?       ���z"@�       �                   ��?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?�       �                  �(S?      �<       z�5��@������������������������       �               ��#�� @������������������������       �               ��#��@������������������������       �               ���>��@�       �                  �6��?v%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?�       �                 �/��?Bǵ3���?       �q�ͨ�@������������������������       �               �cp>@�       �                ��#+y?��Z�	7�?       j~���@�       �                 @�w�?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               ��#���?�       �                 x��?������?       �4^$4�#@�       �                  ��?      �<       �cp>@������������������������       �               ��/����?������������������������       �               0����/@�       �                  0Y��?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@�       �                �o|?~y��]0�?       ���y"@������������������������       �               ��+��+@������������������������       �      ȼ       ��/����?�       �                  {�?BC��?       �WDl��0@�       �                 @L۝?$ k�Lj�?       �q��l}#@�       �                  �k�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ��       ���-��@�       �                 ��=�?���1p8�?       |곯�@������������������������       �               ��#���?�       �                 `TQ�?|��`p��?       �����@������������������������       �               H�4H�4@�       �                 �$��?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?�       �                 ХJ�?%O�f�?       �Q�K�?@�       �                 ��h�?���b�?       �{u;y�-@�       �                �'F�s?$ k�Lj�?       �q��l}@������������������������       �      ��       �cp>@�       �                 ��J�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��+��+$@�       �                  �P�?d�Ѿ�?       ޓr�0@������������������������       �               ��#�� @�       �                  0�9�?x9����?
       }��.�,@�       �                 �8%�?@��~d��?	       8E���*@�       �                 ��Ƚ?���mf�?       毠�?b@������������������������       �               0#0#�?������������������������       �      �<       ��/���@�       �                   �?      �<       E�JԮD!@������������������������       �               ��/����?������������������������       �               ��/���@������������������������       �               0#0#�?�       �                 p�sE?����|e�?       �L���3@������������������������       �               #0#0&@�       �                 ���?�����?       �v�qp�!@������������������������       �               0����/@������������������������       �               0#0#@�       �                 p�:�?���9�۵?%       N}d	�P@�       �                 �E�?d����?       �����!@������������������������       �      ��       �C=�C=@������������������������       �      �<       ��/����?�       �                  �E�? ���:k�?       +��ߵK@�       �                 ���?�^�F�M�?       ��ޚ�&@�       �                 m���?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               vb'vb'"@������������������������       �      ��       #0#0F@�t�bh�hhK ��h��R�(KK�KK��h �B8  �5��P>b@Y���d@�6k�6�c@�,����W@����\@����M@f:��,&S@��/���N@H�4H�4@��#�� @�cp>@        ��#�� @                        �cp>@                ��/����?                ��/���@        �k(��R@�a#6�K@H�4H�4@"�}��P@��|��<@H�4H�4@�P^Cy?@0����/@        ��#���?��/���@        ��#���?                        ��/���@        Kp�}>@��/����?        �#���9@                ��#��@��/����?        ��#��@                        ��/����?        �YLg1B@�e�_��7@H�4H�4@��#��@��On�(@0#0#�?z�5��@                ��#���?��On�(@0#0#�?��#���?鰑%@        ��#���?��/����?                ��/����?        ��#���?                        0����/#@                ��/����?0#0#�?        ��/����?                        0#0#�?���b:@@�cp>'@0#0# @��#�� @���-��@0#0# @z�5��@��/����?        ��#��@                ��#�� @��/����?                ��/����?        ��#�� @                ��#�� @�cp>@0#0# @        �cp>@        ��#�� @        0#0# @��#�� @                                0#0# @�,����7@0����/@        ��#�� @�cp>@        ��#�� @                        �cp>@        �k(���5@��/����?        ��#�� @��/����?        ���>��@                ��#���?��/����?        ��#���?                        ��/����?        ��b:��*@                ��#���?                {�5��(@                ���>��@���-��:@H�4H�4@z�5��@���-��:@0#0#�?z�5��@���-��:@        ��#�� @�cp>�9@        ��#���?�cp>7@                D�JԮD1@        ��#���?�cp>@                �cp>@        ��#���?�cp>@        ��#���?                        �cp>@                ��/����?                ��/����?        ��#���?�cp>@        ��#���?                        �cp>@        ��#���?��/����?                ��/����?        ��#���?                                0#0#�?��#��@        0#0# @��#���?        0#0# @                0#0# @��#���?                z�5��@                �k(��2@n��F:lI@������J@�k(��2@��On�H@�;�;;@�k(��2@	�cp>G@0#0#0@�k(��2@/����/3@#0#0&@ZLg1��&@9l��F:2@0#0#@�k(��"@��/����?0#0# @                0#0# @�k(��"@��/����?        ��#��@��/����?        ��#��@                        ��/����?        ;��,��@                ��#�� @                z�5��@                ��#�� @D�JԮD1@0#0# @��#���?D�JԮD1@        ��#���?���-��@                0����/@        ��#���?��/����?        ��#���?                        ��/����?                鰑%@        ��#���?        0#0# @                0#0# @��#���?                ���>��@��/����?�C=�C=@���>��@��/����?0#0#@                H�4H�4@���>��@��/����?0#0#�?;��,��@                ��#�� @��/����?0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?��#�� @                                H�4H�4@        ���-��:@��+��+@        ��/����?H�4H�4@        ��/����?                        H�4H�4@        �cp>�9@0#0# @        �cp>�9@0#0#�?        ��On�8@                ��/����?0#0#�?                0#0#�?        ��/����?                        0#0#�?        ��/���@#0#0&@        ��/���@0#0#�?                0#0#�?        ��/���@                        ��+��+$@        ��/����?��8��8:@                #0#06@        ��/����?0#0#@        ��/����?0#0#�?        ��/����?                        0#0#�?                H�4H�4@�}�\I@���-��J@f'vb'�X@�}�\I@o��F:lI@��)��)C@�}�\I@	�cp>G@%S2%S27@�,����G@�_��e�=@#0#0&@�GpAF@%jW�v%4@�C=�C=@�GpAF@0����/3@0#0# @��#�� @0����/@        ��#�� @                        0����/@        ���#8E@��|��,@0#0# @�P^Cy/@        0#0# @z�5��@        0#0# @z�5��@                                0#0# @�k(��"@                ��b:��:@��|��,@        ��#��@                \Lg1��6@��|��,@        ������3@��/���@        ��#��0@�cp>@        �P^Cy/@��/����?        ��#�� @��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        z�5��@                ��#�� @                ��#��@                ���>��@                ��#���?��/����?                ��/����?        ��#���?                z�5��@0����/@                �cp>@        z�5��@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ��#���?                z�5��@���-��@                �cp>@                ��/����?                0����/@        z�5��@��/����?                ��/����?        z�5��@                        ��/����?��+��+@                ��+��+@        ��/����?        z�5��@0����/#@0#0#@��#�� @��/���@        ��#�� @��/����?                ��/����?        ��#�� @                        ���-��@        ��#���?��/����?0#0#@��#���?                        ��/����?0#0#@                H�4H�4@        ��/����?0#0#�?        ��/����?                        0#0#�?z�5��@On��O0@H�4H�4(@��#���?��/���@��+��+$@��#���?��/���@                �cp>@        ��#���?��/����?                ��/����?        ��#���?                                ��+��+$@��#�� @��On�(@0#0# @��#�� @                        ��On�(@0#0# @        ��On�(@0#0#�?        ��/���@0#0#�?                0#0#�?        ��/���@                E�JԮD!@                ��/����?                ��/���@                        0#0#�?        0����/@�A�A.@                #0#0&@        0����/@0#0#@        0����/@                        0#0#@        �cp>@+��+��N@        ��/����?�C=�C=@                �C=�C=@        ��/����?                ��/����?�;�;K@        ��/����?��+��+$@        ��/����?0#0#�?        ��/����?                        0#0#�?                vb'vb'"@                #0#0F@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ"�a,hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKم�h��Bx/         �                 0�0�?$��^UT�?,      �	[|�}@                        ���b?��D���?�       I%᎝�s@       p                  �{��?��Y'Ib�?�       m��W��q@       Q                 ��@�?1�嶏�?�       7H�4HCp@       P                 �a�?��:4��?z       �l���ig@       9                 P^N<?���$�?w       hy��f@                        ��u?��3E�?S       ������_@                         .:q?���cE��?4       d�coU@	                        ЮU?V*�"�?0       hܤ?[�S@
                        N��S?�^�#΀�?       O�{��A%@                         �u��?)���?       y��uk!@������������������������       �               ��#���?������������������������       �               ��/���@������������������������       �               ��/����?                        `D*a?t���X��?)       �f�� �P@                        @Ws�?l�s�	�?(       "ߌ��P@                        0��?�<켴��?       �����E@                        �j�%?$Bms�?       ��֖��;@������������������������       �               z�5��(@                        �*f�?M�����?
       p����.@������������������������       �      �<       {�5��(@                        P�W?^%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?                        ,*����B���?	       F��,�,@������������������������       �               �cp>@������������������������       �               [Lg1��&@������������������������       �               |�5��8@������������������������       �      	�       ��/����?������������������������       �               ���>��@       4                 �j�?i;�\q�?       E�c�eD@        %                 pA}?n���;��?       �ڴ���B@!       $                 0��?& k�Lj�?       �q��l}#@"       #                 �؉�?)���?       y��uk!@������������������������       �               ��#���?������������������������       �               ��/���@������������������������       �      ܼ       ��#���?&       +                 �{��?�)z� ��?       ��\�<@'       *                   +Y�?��I@�?       �2d�%@(       )                 �C8�?$ k�Lj�?       �q��l}#@������������������������       �               ��#�� @������������������������       �      ��       ��/���@������������������������       �      ܼ       ��#���?,       3                 �Oc�?j����?       $c�Z%K1@-       0                   \��?bn����?
       � ��w<(@.       /                  'V�?\����?       P	K��@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?1       2                 hՖ�?4=�%�?       �(J��@������������������������       �               ��#�� @������������������������       �               �cp>@������������������������       �               ;��,��@5       6                 �/��?~��`p��?       �����@������������������������       �               0#0#�?7       8                 ���?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?:       E                 ��H?X�ђ���?$       g���J@;       <                 �u)�>��|��?       ó�̙4@������������������������       �               ��#�� @=       B                 @��?�FS�5�?       ��9Շ2@>       ?                 0�aD?�d��}�?       ��Se+@������������������������       �      ��       鰑%@@       A                 @S��?j%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?C       D                  ���?�Z�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@F       I                  s��?�h��%�?       �1�
�u@@G       H                  ;��?      �<       鰑5@������������������������       �               ��/����?������������������������       �               1����/3@J       O                 �(co?b%@�"�?       ��[�'@K       L                 �$I�?���/��?       V��7�@������������������������       �               ��/����?M       N                 ׯ?`n����?       � ��w<@������������������������       �               ��#��@������������������������       �      �<       ��/����?������������������������       �               ��/���@������������������������       �               ���>��@R       g                 |�L?�%�!��?)       �G�:R@S       `                 0p�:?��r�Kk�?       .GnΏ�G@T       U                  �Q�?�i�0��?       ;����?@������������������������       �        
       �C=�C=,@V       _                  P���?�S�p��?	       Q���1@W       \                    �?��;�B(�?       ����*(@X       [                 `0��?���WW�?       �j�S@Y       Z                  �3��?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      �<       z�5��@]       ^                   .p�?Hy��]0�?       ���y"@������������������������       �               ��/����?������������������������       �               ��+��+@������������������������       �               �cp>@a       f                 `�~�?RG�u�?
       ALx��.@b       e                 �3e�?��&���?	       ��G2��,@c       d                 �j��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��On�(@������������������������       �               0#0#�?h       i                  @mj�?&|�!f�?       )�\S'y9@������������������������       �               �cp>'@j       o                 �'��?���/��?       J9U6�+@k       n                 ��ݭ?@���'0�?       �C�� T"@l       m                 �I�w?      �<       ���>��@������������������������       �               z�5��@������������������������       �               ��#��@������������������������       �      �<       ��/����?������������������������       �               0����/@q       |                 ����?�;��sJ�?       ���5�F6@r       w                  <��?�����?       ��ȋ_)2@s       t                 (�Q�?�d�$���?       �T�f@������������������������       �               z�5��@u       v                  ��{�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?x       {                 ���?�n���k�?       3��&�*@y       z                 `z\�?|��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               ��+��+$@}       ~                 PƷ�?�zœ���?       IG���t@������������������������       �               z�5��@������������������������       �               0#0#�?�       �                 0���?�In�� �?       �+�i�@@�       �                  �JV�?w�;B��?       ֟���	@@������������������������       �               �cp>@�       �                  `���?H����D�?       ���2=@�       �                 ����?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               ��8��8:@������������������������       �      �<       ��/����?�       �                 ��5�?�А�X��?f       �#Q��uc@�       �                 0vb�?�B��2�??       � �~g�W@�       �                 ��>�?��4'�?       ~U����C@�       �                 p)j�?���xg��?       �z�+@�       �                 �mx�?��3Fi�?       :�"Ξs@������������������������       �               ��#�� @������������������������       �               ��+��+@�       �                    �?��n��?       �-H�\@�       �                 0���?��q�R�?       C}Ԥ@������������������������       �               ��#���?�       �                  �0��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       ��/���@�       �                 ��Ҧ?�g���E�?       �m���9@������������������������       �      м       0#0#0@�       �                 l��?��G���?       �֔�Э#@�       �                 8���?��[����?       Hl�_A@������������������������       �               0����/@������������������������       �               0#0# @������������������������       �               H�4H�4@�       �                 p&��?�t�� ��?%       ��4�WK@�       �                 Pzo�?Ă����?       K�䙶8@�       �                 p
��?�(1k��?       �ꁞ9�6@�       �                  �E�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @�       �                 �~��?      �<       ������3@������������������������       �               ��#�� @������������������������       �               ��,���1@������������������������       �               0#0# @�       �                 p��?Bʁ���?       ����=@�       �                 �o��?�`Y>�?       Qm�ӽ 6@�       �                  ���?�g�vw�?       {q�^*2@�       �                 P���?�a����?	       AC6&@�       �                 ���?|�G���?       ��%�|@������������������������       �               ��/����?�       �                 ��W�?|��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?�       �                  �?d����?       P	K��@������������������������       �               ;��,��@�       �                 ��y�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               �C=�C=@�       �                 �c�c?      �<       ��/���@������������������������       �               �cp>@������������������������       �               ��/����?�       �                  `�J�?����|e�?       �z �B�@�       �                 6u�?`�ih�<�?       ��
@�       �                 H9A�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��+��+@������������������������       �      ȼ       ��/����?�       �                   ��?�t�yHw�?'       ,N�c'�N@�       �                   �P�?k<S>	�?       T܃���4@�       �                 @Q�?�Rn*l�?       5���2@�       �                 p�͢?r�C7�?       ���7��)@�       �                 �4�?     ��?       "F�b@������������������������       �               ��#�� @������������������������       �               H�4H�4@�       �                 xb'�?pLU���?       i�ҹ^�@������������������������       �               ���-��@������������������������       �               0#0#�?������������������������       �               H�4H�4@������������������������       �      �<       ��#�� @�       �                 @���?�Z}��K�?       `��D@�       �                 �8U|?����/�?       ��
C@�       �                 �L��?p�~:��?       �����)@������������������������       �               0#0#@�       �                 �;�?�����?       �v�qp�!@�       �                 p*�?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �      ��       0����/@������������������������       �               H�4H�4@������������������������       �      ��       k�6k�69@�       �                 H�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?�t�bh�hhK ��h��R�(KK�KK��h �BX  ��k(/d@�z����c@�؉��Ic@	�#�O_@����/k_@:��8�cP@	�#�O_@y�����]@�z��z�B@    �]@�����]@H�4H�48@{�YL�Z@������S@0#0# @�5��X@������S@0#0# @�GpAV@����z�A@0#0# @��,���Q@��/���.@        &�}��O@��/���.@        ��#���?/����/#@        ��#���?��/���@        ��#���?                        ��/���@                ��/����?        �P^CyO@�cp>@        �P^CyO@0����/@        �k(��B@0����/@        �#���9@��/����?        z�5��(@                ��b:��*@��/����?        {�5��(@                ��#���?��/����?                ��/����?        ��#���?                ZLg1��&@�cp>@                �cp>@        [Lg1��&@                |�5��8@                        ��/����?        ���>��@                �k(��2@&jW�v%4@0#0# @�k(��2@/����/3@        ��#�� @��/���@        ��#���?��/���@        ��#���?                        ��/���@        ��#���?                ��#��0@�cp>'@        z�5��@��/���@        ��#�� @��/���@        ��#�� @                        ��/���@        ��#���?                ��b:��*@��/���@        ��#�� @��/���@        z�5��@��/����?        z�5��@                        ��/����?        ��#�� @�cp>@        ��#�� @                        �cp>@        ;��,��@                        ��/����?0#0# @                0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?        <��,��$@��]�ڕE@        z�5��@��|��,@        ��#�� @                ��#��@��|��,@        ��#���?��On�(@                鰑%@        ��#���?��/����?                ��/����?        ��#���?                z�5��@��/����?                ��/����?        z�5��@                ��#��@��|��<@                鰑5@                ��/����?                1����/3@        ��#��@��/���@        ��#��@��/���@                ��/����?        ��#��@��/����?        ��#��@                        ��/����?                ��/���@        ���>��@                [Lg1��&@������C@#0#06@��#��@鰑5@#0#06@z�5��@��/���@��-��-5@                �C=�C=,@z�5��@��/���@�C=�C=@z�5��@��/����?�C=�C=@z�5��@��/����?0#0# @        ��/����?0#0# @        ��/����?                        0#0# @z�5��@                        ��/����?��+��+@        ��/����?                        ��+��+@        �cp>@        ��#���?���-��*@0#0#�?��#���?���-��*@        ��#���?��/����?                ��/����?        ��#���?                        ��On�(@                        0#0#�?���>��@;l��F:2@                �cp>'@        ���>��@���-��@        ���>��@��/����?        ���>��@                z�5��@                ��#��@                        ��/����?                0����/@        ���>��@��/����?��8��8*@��#��@��/����?H�4H�4(@��#��@��/����?        z�5��@                ��#���?��/����?                ��/����?        ��#���?                        ��/����?H�4H�4(@        ��/����?0#0# @                0#0# @        ��/����?                        ��+��+$@z�5��@        0#0#�?z�5��@                                0#0#�?        �cp>@�C=�C=<@        ��/���@�C=�C=<@        �cp>@                ��/����?�C=�C=<@        ��/����?0#0# @        ��/����?                        0#0# @                ��8��8:@        ��/����?        �YLg1B@��/���>@#0#0V@�P^Cy?@0����/3@#0#0F@z�5��@0����/#@�;�;;@z�5��@0����/@H�4H�4@��#�� @        ��+��+@��#�� @                                ��+��+@��#���?0����/@0#0#�?��#���?��/����?0#0#�?��#���?                        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/���@                0����/@��-��-5@                0#0#0@        0����/@��+��+@        0����/@0#0# @        0����/@                        0#0# @                H�4H�4@,�����;@0����/#@S2%S2%1@�k(���5@��/����?0#0# @�k(���5@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ������3@                ��#�� @                ��,���1@                                0#0# @z�5��@D�JԮD!@�A�A.@z�5��@���-��@vb'vb'"@z�5��@�cp>@vb'vb'"@z�5��@�cp>@0#0# @        ��/����?0#0# @        ��/����?                ��/����?0#0# @                0#0# @        ��/����?        z�5��@��/����?        ;��,��@                ��#���?��/����?                ��/����?        ��#���?                                �C=�C=@        ��/���@                �cp>@                ��/����?                ��/����?H�4H�4@        ��/����?H�4H�4@        ��/����?0#0#�?        ��/����?                        0#0#�?                ��+��+@        ��/����?        ;��,��@�cp>'@#0#0F@��#��@���-��@��+��+$@��#�� @���-��@��+��+$@��#�� @���-��@0#0#@��#�� @        H�4H�4@��#�� @                                H�4H�4@        ���-��@0#0#�?        ���-��@                        0#0#�?                H�4H�4@��#�� @                ��#���?0����/@T2%S2%A@        0����/@B�A�@@        0����/@0#0# @                0#0#@        0����/@0#0#@        0����/@0#0#�?                0#0#�?        0����/@                        H�4H�4@                k�6k�69@��#���?        0#0#�?��#���?                                0#0#�?�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�8�hhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK���h��B6         �                 ���b?6�z�tL�?2      ����u�}@       �                 �'>�?��D�|��?�       ���.w@       �                 ��U�?;[���?�       �"��u@       a                 �Շ�?r��	�r�?�       {)G_p@                        �`>R?�q�)r�?p       �#zef@                        P�_?^dؗ��?       4d��8@                        0��>�)z� ��?       ��\�@       	                 `���>Δfm���?       ��Z�N@������������������������       �               ��#���?
                        � ^P?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               z�5��@                         �u��?v@ȱ��?       ���~1@������������������������       �               ��#���?                        �
;E?�h��%�?
       �1�
�u0@                        j��Q?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      ��       ���-��*@       T                 @�:�?�D��?a       �57Uc@       ;                 )DW?���8j��?O       #��h�]@       :                 �x{}?L��Z%�?3       ��V&b�R@       #                   �G�?��e����?1       J';d�Q@       "                    �?��R ��?	       ⲿꁞ+@                         �#n?>9�)\e�?       _���b @������������������������       �               ��/����?       !                 pZW?�����?       �O��@                         Pmj�?bn����?       � ��w<@������������������������       �               ��#���?                          `�J�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               z�5��@������������������������       �      ȼ       �cp>@$       9                 P�ba?X�־+��?(       �I��'3L@%       6                  ���?�s���?       [E��K�C@&       3                 (߁C?H1`f+q�?       6�W���?@'       0                 r�4?h�j���?       ^��\�;@(       -                 �\͵?���Ѯ�?
       ��GQ&@)       *                 8�,�?��6L�n�?       �E#��h @������������������������       �      �<       z�5��@+       ,                 ��aӾ���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?.       /                  `���?V%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?1       2                  �.�?      �<       ��#��0@������������������������       �               ��#�� @������������������������       �               ���>��,@4       5                    �?      �<       ��/���@������������������������       �               ��/����?������������������������       �               ��/����?7       8                    �?      �<       ��#�� @������������������������       �               ���>��@������������������������       �               ��#���?������������������������       �        	       ��#��0@������������������������       �               0����/@<       O                 0I��?|�+�ޯ�?       V4�@�E@=       H                 @���?�Ug���?       ����@@>       E                  ���?��/ʪ��?       I�Ų��1@?       D                 �U�,?�F���?       :�.�-'@@       A                 ��Y?`�r{��?       e�6� @������������������������       �               ��/���@B       C                  oEg?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               ��/���@F       G                 Hl�f?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#��@I       N                   ���?TF�X��?	       .�=k�U0@J       K                  %�r?M�����?       p����.@������������������������       �               [Lg1��&@L       M                 @�r�?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      м       ��/����?P       Q                  ����?ܜ�x�?       d��إV#@������������������������       �               0����/@R       S                 `�h'?  k�Lj�?       �q��l}@������������������������       �               ��#���?������������������������       �      �<       ��/���@U       X                  p��?��k\��?       nG�
 B@V       W                 8�{?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @Y       Z                 �'�?�C=+��?       c��T|@@������������������������       �               ��/����?[       `                 �	�}?�)��ĭ?       ��[��@@\       ]                 hI�P?�FO���?       �ߌ$@������������������������       �               ��#�� @^       _                 ��[?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �        	       �k(���5@b       g                 �\�?�4 ��?1       ���\(�T@c       f                  L��?�}	;	�?       vK�>4%@d       e                 x��?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?������������������������       �               ��/���@h       �                 0�{?4" PD��?,       K:�}�R@i       n                   ��?��g��B�?       ����;B@j       m                 0}}?�^�#΀�?       O�{��A%@k       l                 p��!?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      �<       ��/���@o       z                 @�r�?�x��>�?       �	�{ �9@p       y                 ��Z�? $�W �?	       �xy'�)@q       x                 �H�y?�Wf]�?       ?���g�!@r       s                    �?��d
���?       f�G�N�@������������������������       �               �cp>@t       u                 ��d?b,���O�?       ���/>@������������������������       �               0#0# @v       w                  #3x?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               0#0# @������������������������       �      ��       ��/���@{       �                  ��d�?$��C/��?       �~*@|       }                 �6��?D��NV=�?       �t�ܲ@������������������������       �               ��/����?~                         @V��?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               vb'vb'"@�       �                 `�e�?�8u#��?       ��_O;�A@�       �                 �$�?!��8���?       �<z z*@������������������������       �               z�5��@�       �                 p� �?��[����?       Hl�_A@������������������������       �               0#0# @������������������������       �               0����/@�       �                 ��m�?�(1k��?       �ꁞ9�6@�       �                 ����?\����?       P	K��@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?������������������������       �      �<       �P^Cy/@�       �                 �*��?�)���?;       p�m�U3U@�       �                  ��?�2+xa��?       �|�hrE4@�       �                    �?�O
�*Q�?       �͉V�M2@�       �                 `�A�?$ k�Lj�?       �q��l}@������������������������       �      ��       �cp>@�       �                  ���?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 �\͵?      �<	       ���-��*@������������������������       �               ��/����?������������������������       �               �cp>'@�       �                 �s��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 p5W�?��*���?+       4K4
�!P@�       �                 <�Q?��5��`�?#       '�1��H@�       �                 ���?06����?       �OY�9D@�       �                 �%��?d�����?       N��P�B@�       �                  �?�Z�ѕ�?       ��G3l?@�       �                 �=M�?����h�?       @��o{3@�       �                  `S��?��^���?       ���w1@�       �                 @Ws�?.�8�4�?       ׁ��t0@�       �                   .p�?z�G���?       '5L�`�@������������������������       �               0#0# @�       �                 ��`�?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �        	       鰑%@������������������������       �               0#0#�?������������������������       �               0#0# @�       �                 @咣?���R�?       f��R�'@������������������������       �               ;��,��@�       �                 @� ?�;�a
=�?       ��l��@������������������������       �               ��/���@�       �                 �{��?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 ��?�y��]0�?       ���y"@������������������������       �               ��/����?������������������������       �               ��+��+@������������������������       �      �       H�4H�4@�       �                 ���?��r{��?       e�6� @������������������������       �               ��/���@�       �                 ����?Ɣfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@�       �                 `���?�W���?       �4m��T0@�       �                 @��8?�/,Tg�?       �����*@�       �                 �@�?     ��?       "F�b@������������������������       �               ��#�� @������������������������       �               H�4H�4@������������������������       �               ��#�� @�       �                �g�?j%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 h��?4��
�t�?       �r�%6@�       �                  ;��?`�ih�<�?       W�3D*5@�       �                �\�ѓ?|��`p��?       �����@������������������������       �               0#0#�?�       �                 (H?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 �P�?d*�'=P�?        �22@������������������������       �               ��/����?�       �                 �$I�?�6��b�?
       &�|�1@������������������������       �               ��8��8*@�       �                 p4N�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �      �<       ��#���?�       �                 @4��?�n<��i�?G       �Cc��Y@�       �                 ��<{?�������?0       "�WQ@������������������������       �               ��#���?�       �                 ��|�?�Q�X��?/       �T�tQ@�       �                  �ni?��#���?       �͆�1�2@������������������������       �               ��/����?�       �                 0#ή?��i���?       ����1@�       �                 �YJ�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                 �.K�?�n���k�?
       3��&�*@�       �                 ��a�?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?������������������������       �               0#0# @�       �                 8�C�?@-�0���?"       �B�?O�H@������������������������       �               dJ�dJ�A@�       �                  N��?P��ճC�?       y��l$,@������������������������       �        	       H�4H�4(@�       �                 ����?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 `j��?xT`�[k�?       �m����@@�       �                 ��~?P�b��?       ���"7@������������������������       �               ��/����?�       �                  ��?�~���9�?       �q�Ί#6@�       �                  Y��?Hy��]0�?       ���y"@�       �                 �M�?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      ��       H�4H�4@������������������������       �        
       0#0#0@�       �                 �)��?(�Jg@��?       ��G� �%@�       �                 ��*�?�;�a
=�?       ��l��@������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �               0#0#@�t�bh�hhK ��h��R�(KK�KK��h �B(  Qg1���d@F:l��d@xb'vb'b@?��,��d@��z��wb@�+��+�K@-�����d@W<�œb@�z��z�B@�5��P>b@t%jW�vX@vb'vb'2@��P^C�\@��P@        ���>��@E�JԮD1@        ��#��@�cp>@        ��#���?�cp>@        ��#���?                        �cp>@                ��/����?                ��/����?        z�5��@                z�5��@��|��,@        ��#���?                ��#�� @��|��,@        ��#�� @��/����?        ��#�� @                        ��/����?                ���-��*@        ��b:��Z@��h
�G@        �k(��R@h
��F@        �>��nK@%jW�v%4@        �>��nK@��/���.@        ;��,��@E�JԮD!@        ;��,��@�cp>@                ��/����?        ;��,��@��/����?        ��#�� @��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                z�5��@                        �cp>@        ~�5��H@���-��@        ��#��@@���-��@        }�5��8@���-��@        |�5��8@�cp>@        ��#�� @�cp>@        ���>��@��/����?        z�5��@                ��#���?��/����?                ��/����?        ��#���?                ��#���?��/����?                ��/����?        ��#���?                ��#��0@                ��#�� @                ���>��,@                        ��/���@                ��/����?                ��/����?        ��#�� @                ���>��@                ��#���?                ��#��0@                        0����/@        ������3@�e�_��7@        �k(��2@��/���.@        ;��,��@��On�(@        ��#���?鰑%@        ��#���?���-��@                ��/���@        ��#���?�cp>@        ��#���?                        �cp>@                ��/���@        ��#��@��/����?                ��/����?        ��#��@                ��b:��*@�cp>@        ��b:��*@��/����?        [Lg1��&@                ��#�� @��/����?        ��#�� @                        ��/����?                ��/����?        ��#���?E�JԮD!@                0����/@        ��#���?��/���@        ��#���?                        ��/���@        ��#��@@�cp>@        ��#�� @��/����?                ��/����?        ��#�� @                �P^Cy?@��/����?                ��/����?        �P^Cy?@��/����?        �k(��"@��/����?        ��#�� @                ��#���?��/����?                ��/����?        ��#���?                �k(���5@                �P^Cy?@�-����@@vb'vb'2@        0����/#@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/���@        �P^Cy?@�e�_��7@S2%S2%1@z�5��@9l��F:2@�A�A.@��#���?/����/#@        ��#���?��/����?        ��#���?                        ��/����?                ��/���@        ��#�� @D�JԮD!@�A�A.@��#���?���-��@��+��+@��#���?�cp>@��+��+@��#���?�cp>@H�4H�4@        �cp>@        ��#���?        H�4H�4@                0#0# @��#���?        0#0#�?��#���?                                0#0#�?                0#0# @        ��/���@        ��#���?��/����?��+��+$@��#���?��/����?0#0#�?        ��/����?        ��#���?        0#0#�?                0#0#�?��#���?                                vb'vb'"@*�����;@�cp>@0#0# @z�5��@0����/@0#0# @z�5��@                        0����/@0#0# @                0#0# @        0����/@        �k(���5@��/����?        z�5��@��/����?        z�5��@                        ��/����?        �P^Cy/@                �k(��2@��h
�G@��)��)3@��#���?9l��F:2@0#0#�?��#���?D�JԮD1@        ��#���?��/���@                �cp>@        ��#���?��/����?        ��#���?                        ��/����?                ���-��*@                ��/����?                �cp>'@                ��/����?0#0#�?        ��/����?                        0#0#�?��,���1@��|��<@vb'vb'2@z�5��@���-��:@�A�A.@;��,��@%jW�v%4@�A�A.@;��,��@%jW�v%4@H�4H�4(@;��,��@/����/3@�C=�C=@        ���-��*@H�4H�4@        ���-��*@0#0#@        ���-��*@H�4H�4@        �cp>@H�4H�4@                0#0# @        �cp>@0#0#�?        �cp>@                        0#0#�?        鰑%@                        0#0#�?                0#0# @;��,��@�cp>@0#0#�?;��,��@                        �cp>@0#0#�?        ��/���@                ��/����?0#0#�?                0#0#�?        ��/����?                ��/����?��+��+@        ��/����?                        ��+��+@                H�4H�4@��#���?���-��@                ��/���@        ��#���?�cp>@        ��#���?                        �cp>@        [Lg1��&@��/����?H�4H�4@<��,��$@        H�4H�4@��#�� @        H�4H�4@��#�� @                                H�4H�4@��#�� @                ��#���?��/����?        ��#���?                        ��/����?        ��#���?�cp>@vb'vb'2@        �cp>@vb'vb'2@        ��/����?0#0# @                0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                ��/����?0#0#0@        ��/����?                ��/����?0#0#0@                ��8��8*@        ��/����?H�4H�4@        ��/����?                        H�4H�4@��#���?                ��#���?��On�(@��
�pV@��#���?0����/@T��N��O@��#���?                        0����/@R��N��O@        ��/���@�A�A.@        ��/����?                ��/����?�A�A.@        ��/����?H�4H�4@        ��/����?                        H�4H�4@        ��/����?H�4H�4(@        ��/����?0#0#@                0#0#@        ��/����?                        0#0# @        ��/����?L�4H�4H@                dJ�dJ�A@        ��/����?��8��8*@                H�4H�4(@        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/���@��8��8:@        ��/����?��-��-5@        ��/����?                ��/����?��-��-5@        ��/����?��+��+@        ��/����?0#0# @        ��/����?                        0#0# @                H�4H�4@                0#0#0@        �cp>@��+��+@        �cp>@0#0#�?                0#0#�?        �cp>@                        0#0#@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJP�dhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKυ�h��BH-         �                 �6Sz?��C��S�?2      |��M�z}@       �                 P7&E?n���?�       ��b��w@       z                 �U���ҝu�O��?�       ��I�Xr@       q                 @���?�:%'��?�       L�qBh@       d                 p��?X���?r       |���~e@       [                 @��?��uD�	�?b       ����� b@       :                    �?p���W�?P       �na��2^@                        ���>�ot��?.       Quh�0Q@	                         �Q�?$ k�Lj�?       �q��l}@
                        �;�N?Ɣfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               ��/����?       %                   ��?B��E��?+       41?�O@       "                 �I?��N�?       UQ�dA@                        0�2�?l]ү�8�?       
u-��o8@                         ;��?����ӱ�?       � sE�.0@                        0��?��6L�n�?       �E#��h @                        �i�?����?       ��X�)B@������������������������       �      ��       z�5��@������������������������       �      �<       ��/����?                        Їq?      �<       ��#��@������������������������       �               ��#�� @������������������������       �               ��#�� @                         @?��?���/��?       T��7�@                         ����?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �      м       ��/����?                        �(�?|�t1u�?       "�te!� @������������������������       �               ;��,��@        !                 `0��?N����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @#       $                 0��?      �<       <��,��$@������������������������       �               ��#���?������������������������       �               �k(��"@&       +                 pe�S?�0zQ6W�?       c-�S�=@'       (                 ��?jQ��?       �s�=�!@������������������������       �               0����/@)       *                �3�.s?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @,       7                 NK�X?Ld���?       ��õQ4@-       0                  �Ԧ�?*�q��?       �Mc�(@.       /                  ��d�?b,���O�?       ���/>@������������������������       �               ��#���?������������������������       �               H�4H�4@1       6                 �h�?���/��?       U��7�@2       3                ���`s?�d�$���?       �T�f@������������������������       �               z�5��@4       5                 ��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               �cp>@8       9                 Ȭ�?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ���>��@;       R                 0vb�?&Ϻ���?"       �;���J@<       Q                 @��?$�����?       џ��<@=       P                 ���?Bb
y�	�?       N/㔐k9@>       M                 ��~?�<=��c�?       0ne��Y7@?       H                 ��gn?"Iz�9��?       ��[5@@       E                  _�
?e��}�?	       ��Se+@A       B                 �C[?$ k�Lj�?       �q��l}@������������������������       �               ��/����?C       D                 `���>`%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?F       G                  �~��?      �<       E�JԮD!@������������������������       �               ��/����?������������������������       �               ��/���@I       L                 H��?���`�?       ��
�Me@J       K                 �@�?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               0����/@N       O                 �?�r?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      �<       ��#�� @������������������������       �      ȼ       z�5��@S       Z                 �b)�?hՏ�m|�?       ��h
�7@T       U                 �vQ?��Z�	7�?       j~���$@������������������������       �               ;��,��@V       Y                  �x��?& k�Lj�?       �q��l}@W       X                  ��g�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �      ��       ��b:��*@\       ]                 �m��?h��mf�?       ��b�:8@������������������������       �               0#0#@^       _                  P�"�?�G�<�J�?       S �24@������������������������       �               鰑%@`       a                 �b'�?�5JH���?	       �MOI#@������������������������       �               ��/���@b       c                 T���?z�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?e       f                 @/��?��X<��?       �K��:@������������������������       �               0#0#@g       h                  ��?Φ�a���?       m����6@������������������������       �               0����/@i       p                    �?��b���?       � X�2@j       m                 p5W�?�����?       X!��&@k       l                 �8�?�.�KQu�?       �K̎@������������������������       �               0#0#@������������������������       �               z�5��@n       o                 GW�d?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               �C=�C=@r       s                  @��?HY�����?       ���o]5@������������������������       �               ��/����?t       u                 ����?������?       �_n��4@������������������������       �               #0#0&@v       w                 ՟�?�Wf]�?       ?���g�!@������������������������       �               ��#���?x       y                 8p=�?�~�&��?       ?�]��@������������������������       �               �cp>@������������������������       �               ��+��+@{       �                 �s?���SE>�?<       (�+��W@|       �                 P�c�?��6L�n�?!       ��4}i�H@}       �                 p�R?��k���?       H+զm7F@~       �                 `?�!?����X��?	       (��֞&@       �                 QU�>      �<       �k(��"@������������������������       �               ��#���?������������������������       �               ��#�� @�       �                    �?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#��@@�       �                 Њ�8?      �<       0����/@������������������������       �               ��/����?������������������������       �               �cp>@�       �                 Pܪ�?��=�g]�?       �K��R�F@�       �                 pTF�?�(���?       x��uk1@������������������������       �      ��       �cp>'@�       �                 �n]�?d%@�"�?       ��[�@������������������������       �      �<       ��/���@������������������������       �               ��#�� @�       �                 p�37? �Fl�R�?       ��޷/�<@�       �                 _5?�Wf]�?       ?���g�!@�       �                �٬Ӌ?wT �+��?       ��>Y��@������������������������       �               �cp>@�       �                 (y�?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               H�4H�4@�       �                    �?�U���?
       ����{�3@�       �                 ��?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@�       �                 �Z�?�%�?       �����.@������������������������       �               ��#�� @�       �                 ��N�?,Lj����?       ���T�@������������������������       �               0#0#�?������������������������       �               z�5��@�       �                 0�"]?�/����?>       8�d,�V@�       �                 @� �?�ȁ��?'       ?v�&N@�       �                 ��7?|�:���?%       }F�7�L@�       �                 p���>`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @�       �                 �U*P?<Ό�߂�?"       s�ʽKK@�       �                 P
��?Ы����?       r��9@������������������������       �               ��|��,@�       �                    �?�>s{Ab�?       aI��n'@�       �                 �>��?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �               0����/@������������������������       �      ��       �cp>@�       �                 @�Q?|�y3.��?       �7|	�<@������������������������       �               ��#���?�       �                 �JI�?���C��?       @W=��;@������������������������       �        	       :l��F:2@�       �                 �^7�?�C>�?       �1�m�!@������������������������       �               ��#�� @�       �                 ��>�?�;�a
=�?       ��l��@������������������������       �               �cp>@������������������������       �               0#0#�?�       �                ��1�?H����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @�       �                  ����?nI3%�d�?       ���G�>@�       �                 `9�`?�
���?
       �O���/@������������������������       �               ��#�� @�       �                 �*|}?�Y�Z�?	       U�S��u+@�       �                 ��E�?�g�vw�?       �Aws}8@�       �                  pS��?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               H�4H�4@������������������������       �               ��/���@�       �                 ���o?�)w�q�?       ��|��-@�       �                 pF�?�^�F�M�?
       ��ޚ�&@������������������������       �               ��/����?������������������������       �        	       ��+��+$@�       �                 H��?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@�       �                 `I9�?p�}n Ӯ?8       H�s��(W@�       �                 ��;�?6hh���?       ~�DXR�)@������������������������       �               ��+��+$@������������������������       �      �<       �cp>@������������������������       �        2       �6k�6�S@�t�b�$     h�hhK ��h��R�(KK�KK��h �Bh  y�YLGc@�B�)Dd@��jc@y�YLGc@f
���c@<��8�cP@������a@�œ[<9X@J�4H�4H@������S@����Q@��-��-E@���khS@��t�HQ@��8��8:@��Gp_R@>��18N@#0#0&@��Gp_R@�)�B�D@H�4H�4@]Lg1��F@0����/3@0#0#@��#���?��/���@        ��#���?�cp>@                �cp>@        ��#���?                        ��/����?        �GpAF@��/���.@0#0#@���>��<@0����/@0#0#�?�k(��2@0����/@0#0#�?ZLg1��&@0����/@        ���>��@��/����?        z�5��@��/����?        z�5��@                        ��/����?        ��#��@                ��#�� @                ��#�� @                ��#��@��/���@        ��#��@��/����?                ��/����?        ��#��@                        ��/����?        ���>��@        0#0#�?;��,��@                ��#�� @        0#0#�?                0#0#�?��#�� @                <��,��$@                ��#���?                �k(��"@                �P^Cy/@鰑%@H�4H�4@��#�� @���-��@                0����/@        ��#�� @��/����?                ��/����?        ��#�� @                ��b:��*@��/���@H�4H�4@;��,��@��/���@H�4H�4@��#���?        H�4H�4@��#���?                                H�4H�4@��#��@��/���@        ��#��@��/����?        z�5��@                ��#���?��/����?        ��#���?                        ��/����?                �cp>@        ��#�� @                ��#���?                ���>��@                +�����;@h
��6@0#0# @��#�� @;l��F:2@0#0# @;��,��@9l��F:2@0#0# @z�5��@:l��F:2@0#0# @��#�� @D�JԮD1@0#0# @��#���?��On�(@        ��#���?��/���@                ��/����?        ��#���?��/����?                ��/����?        ��#���?                        E�JԮD!@                ��/����?                ��/���@        ��#���?0����/@0#0# @��#���?        0#0# @��#���?                                0#0# @        0����/@        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                z�5��@                ������3@��/���@        z�5��@��/���@        ;��,��@                ��#���?��/���@        ��#���?��/����?                ��/����?        ��#���?                        �cp>@        ��b:��*@                        1����/3@��+��+@                0#0#@        0����/3@0#0#�?        鰑%@                D�JԮD!@0#0#�?        ��/���@                ��/����?0#0#�?                0#0#�?        ��/����?        ��#��@��/���@�A�A.@                0#0#@��#��@��/���@#0#0&@        0����/@        ��#��@�cp>@#0#0&@��#��@�cp>@0#0#@z�5��@        0#0#@                0#0#@z�5��@                ��#���?�cp>@        ��#���?                        �cp>@                        �C=�C=@��#���?��/���@0#0#0@        ��/����?        ��#���?�cp>@0#0#0@                #0#0&@��#���?�cp>@��+��+@��#���?                        �cp>@��+��+@        �cp>@                        ��+��+@���b:P@��On�8@H�4H�4@�k(���E@�cp>@        �k(���E@��/����?        <��,��$@��/����?        �k(��"@                ��#���?                ��#�� @                ��#���?��/����?                ��/����?        ��#���?                ��#��@@                        0����/@                ��/����?                �cp>@        ;��,��4@0����/3@H�4H�4@��#�� @��/���.@                �cp>'@        ��#�� @��/���@                ��/���@        ��#�� @                �k(��2@��/���@H�4H�4@��#���?�cp>@��+��+@��#���?�cp>@0#0# @        �cp>@        ��#���?        0#0# @��#���?                                0#0# @                H�4H�4@��,���1@��/����?0#0#�?z�5��@��/����?                ��/����?        z�5��@                ���>��,@        0#0#�?��#�� @                z�5��@        0#0#�?                0#0#�?z�5��@                [Lg1��&@2����-O@S2%S2%1@���>��@��On�H@H�4H�4@;��,��@��On�H@0#0# @��#�� @��/����?                ��/����?        ��#�� @                z�5��@y%jW�vH@0#0# @        ��On�8@0#0#�?        ��|��,@                鰑%@0#0#�?        0����/@0#0#�?                0#0#�?        0����/@                �cp>@        z�5��@�e�_��7@0#0#�?��#���?                ��#�� @�e�_��7@0#0#�?        :l��F:2@        ��#�� @�cp>@0#0#�?��#�� @                        �cp>@0#0#�?        �cp>@                        0#0#�?��#�� @        0#0#�?                0#0#�?��#�� @                ��#��@��On�(@�C=�C=,@��#��@D�JԮD!@H�4H�4@��#�� @                ��#�� @D�JԮD!@H�4H�4@��#�� @��/����?H�4H�4@��#�� @��/����?        ��#�� @                        ��/����?                        H�4H�4@        ��/���@                ��/���@#0#0&@        ��/����?��+��+$@        ��/����?                        ��+��+$@        �cp>@0#0#�?                0#0#�?        �cp>@                �cp>@��
�pV@        �cp>@��+��+$@                ��+��+$@        �cp>@                        �6k�6�S@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�g?BhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK���h��B6         �                 ��{�?C"c�O�?2      �FZ5��}@       i                 0-3�?hޜA�F�?'      �
%��H|@       Z                   B�?VV?�E�?x       �qKL�sg@       U                 ����?��鿕��?l       ����&e@       ,                 @ߠs?Y��mk��?f       :�U�@d@       +                 0*��?�̳9��?9       �OG��2X@       *                 P�h�?��~j�X�?7       *�xr��V@                        �94W?x�{7��?2       Å۬QT@	                         y��?�HU����?$       mgP�.TK@
                        "?b����?       ;��18>@������������������������       �        	       \Lg1��&@                        �{�T?�KĈ�?       y�Zc�2@                          ��?��߭Q��?       �QVl�0@������������������������       �               0����/@                        �\ͥ?���/��?       @z$S��'@                           �?��Z�	7�?       j~���$@������������������������       �               z�5��@������������������������       �      �<       ��/���@������������������������       �      ��       ��/����?������������������������       �      ܼ       ��#�� @                        �΢��&��$C�?       ���+p8@                         ��k?(��c`�?       %��t5)@������������������������       �      �<       �cp>'@������������������������       �      ܼ       ��#���?                        �ȠF?�4��v�?       �Y-"�'@                        �/f?�����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?                           �?      �<       �cp>@������������������������       �               �cp>@������������������������       �               �cp>@        !                  Pmj�?�(߫$��?       1H����:@������������������������       �               ��/����?"       '                  ��d�?tb8�Y�?       GJͰ8@#       $                 `��a?X ����?
       1
C>�5@������������������������       �               ��,���1@%       &                 �؉�?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@(       )                  ���?dn����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               <��,��$@������������������������       �               ;��,��@-       R                 0�?�?���va�?-       %�լNP@.       O                 �!�?%���k��?(       \Y@��M@/       D                  #B�?�V�~��?%       �i��L@0       5                 �8{?��c`��?       ���C@1       2                 x��?e��}�?	       ��Se+@������������������������       �      ��       鰑%@3       4                 ����?j%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?6       A                 �~��?bdؗ��?       4d��8@7       8                  ���?�{k���?       P�_�q6@������������������������       �               ��#���?9       :                    �?R�ђ���?       �oFݜh5@������������������������       �               �cp>'@;       <                 ��{?4=�%�?       �(J��#@������������������������       �               0����/@=       @                 �Y�b?�d�$���?       �T�f@>       ?                 H���?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ��       ��#�� @B       C                  ����?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?E       J                    �?ɣ���c�?
       8oU��2@F       G                 0�,�?�<;�`(�?       ��^�&@������������������������       �               ��#��@H       I                   .p�?�w��d��?       �0���s@������������������������       �               H�4H�4@������������������������       �      �<       ��/���@K       N                 `ΐ�?�_�A�?       炵�e`@L       M                 ����?`%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��#��@P       Q                 �%�?~��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @S       T                 ��ى?�����?       �O��@������������������������       �               ��/����?������������������������       �               ;��,��@V       Y                 �m�?P�h��?       S�D'�@W       X                  ��g�?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @������������������������       �               ��#��@[       h                  @���?����X�?       ����f2@\       g                  rp�?ĵM�-�?	       �\�&�.@]       d                 P�h?H[�Jg�?       X�S0f�*@^       c                ��a�?��b�}�?       ���\�@_       `                  ��g�?���/��?       V��7�@������������������������       �               ��/����?a       b                �|�@!?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               0#0#�?e       f                 �m�?      �<       ��#�� @������������������������       �               ��#�� @������������������������       �               z�5��@������������������������       �               0#0# @������������������������       �               z�5��@j       �                 p��?����#�?�       �Q����p@k       �                 0�"]?09����?l       ���Z�e@l       �                 �/�?�Ģ<��?D       3�5O�\@m       �                 �x?>RgO��?1       ѳ��SCU@n                        �U��>Ҕ����?       P@���hF@o       t                 ���?T;պoL�?       ��Xi<@p       q                 ��}w?�}	;	�?       uK�>4%@������������������������       �               �cp>@r       s                 @Ͻ}?���mf�?       毠�?b@������������������������       �               0#0#�?������������������������       �      �<       ��/���@u       ~                 ��?����?       8��9�1@v       }                  0B�?�}/W�?       �r�.�%@w       |                  Џ~�?z�G���?       ��%�|@x       {                   E(�?���mf�?       毠�?b@y       z                  ����?~�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �               H�4H�4@������������������������       �               �cp>@������������������������       �               �C=�C=@�       �                 ���f?ॏje��?	       ��BLGh0@������������������������       �               0#0# @������������������������       �               ��|��,@�       �                  �g<�?�݄s�w�?       W'�$�D@�       �                  y��?v@ȱ��?       om���S'@�       �                 @?      �<       D�JԮD!@������������������������       �               ��/����?������������������������       �               ���-��@�       �                 @���?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?�       �                 ��7�?��Q���?       ��Ǒ<@�       �                 P=)�?`��qS�?       �X���0@�       �                  ��>�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �        	       ���>��,@�       �                 ��ٹ?�3`���?       �~�M�(@������������������������       �               z�5��@�       �                 p��?|��`p��?       f;3@��!@�       �                 ���?`�ih�<�?       ��
@�       �                  pS��?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?�       �                  ��u�?�!vi��?       �qw1;@�       �                 ��&�?N��L��?       ��G��8@�       �                  s��?PR9�� �?       ���55  @�       �                 �ƽ?�@G���?       hu��@������������������������       �               ��/����?�       �                 (p�J?~�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                ��Sl�?�zœ���?       IG���t@������������������������       �               0#0#�?������������������������       �               z�5��@�       �                 �%��?r����?       Qz�i0@�       �                 �и?X�ih�<�?       ��
@������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?������������������������       �      ��       vb'vb'"@������������������������       �      ȼ       z�5��@�       �                 ��c�?ʒ�0�?(       ��G�O@������������������������       �      ȼ       �
��
�E@�       �                 p@�?�&t�ׁ�?       4�1!�4@�       �                 �%{�?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?�       �                 p1m�?7��b�?       &�|�1@������������������������       �        	       �A�A.@�       �                 v�2�?��G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 �\��?J��Z*:�?C       ~�#�RV@�       �                 �TI�?����K�?       5�(��3@�       �                 py?����U�?       5�ժ�c)@������������������������       �               H�4H�4@�       �                 @��?�ۜ�x�?	       c��إV#@�       �                 P�2<?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �      ��       ���-��@�       �                 x�׀?�AP�9��?       i��6��@������������������������       �               ��/����?������������������������       �               ��+��+@�       �                 �6SZ?�)A��e�?3       �PY�hQ@�       �                 ���?�LgF��?$       Ɖ�E�GI@�       �                  �G?V�wi�*�?"       UK�^v�G@�       �                 p��?ع����?       T6���B@�       �                �s�[w?l����s�?       ��/�StA@�       �                 ��:�?��P����?       ;#��,@ @������������������������       �               ��/����?�       �                   .p�?k��9�?       �J���@������������������������       �               z�5��@�       �                 �Y��?b,���O�?       ���/>@�       �                 �x��?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               0#0# @�       �                  �^��?�F�o��?       (��:@������������������������       �               ��/����?�       �                 P���?�z��o�?       1�����9@������������������������       �               ������3@�       �                 X��?T����1�?       ��;9�@������������������������       �               0#0# @������������������������       �               ��#��@�       �                  �JV�?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?�       �                   ҏ�?"4=�%�?       �(J��#@�       �                 0���?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@�       �                 �m��?r@ȱ��?       om���S@������������������������       �               ��#���?������������������������       �               0����/@�       �                 �5W�?     ��<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?�       �                  ��?H?�	,�?       >0�1b3@������������������������       �               ��+��+$@�       �                    �?d����?       �����!@������������������������       �               H�4H�4@�       �                 Pα�?z��`p��?       �����@�       �                 � ğ?�� ��?       rp� k@������������������������       �               ��/����?�       �                  ���?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               H�4H�4@�       �                 �+�[?��R���?       :�S) 4@�       �                 �-�?     ��?       "F�b@������������������������       �               0#0# @�       �                 �@�?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?�       �                 �t_�?��E�B��?       dߞKC.@������������������������       �               ��/����?������������������������       �               ��8��8*@�t�bh�hhK ��h��R�(KK�KK��h �B(  cCy��d@�+Q��b@��jc@?��,��d@��z��wb@`��[�ea@V^CyeZ@}����Q@��+��+$@���W@M!��Q@�C=�C=@�k(���U@M!��Q@��+��+@���b:P@On��O@@            �M@Pn��O@@        6��tSH@On��O@@        �#���9@��|��<@        ������3@鰑%@        \Lg1��&@                ��#�� @鰑%@        z�5��@鰑%@                0����/@        z�5��@�cp>@        z�5��@��/���@        z�5��@                        ��/���@                ��/����?        ��#�� @                z�5��@:l��F:2@        ��#���?�cp>'@                �cp>'@        ��#���?                ;��,��@���-��@        ;��,��@��/����?        ;��,��@                        ��/����?                �cp>@                �cp>@                �cp>@        [Lg1��6@��/���@                ��/����?        [Lg1��6@��/����?        ;��,��4@��/����?        ��,���1@                z�5��@��/����?                ��/����?        z�5��@                ��#�� @��/����?                ��/����?        ��#�� @                <��,��$@                ;��,��@                \Lg1��6@�+Q��B@��+��+@��,���1@=l��F:B@��+��+@��,���1@����z�A@H�4H�4@��#�� @�_��e�=@        ��#���?��On�(@                鰑%@        ��#���?��/����?        ��#���?                        ��/����?        ���>��@D�JԮD1@        ;��,��@D�JԮD1@        ��#���?                ��#��@D�JԮD1@                �cp>'@        ��#��@�cp>@                0����/@        ��#��@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ��#�� @                ��#�� @                ��#���?                ��#���?                �k(��"@�cp>@H�4H�4@��#��@��/���@H�4H�4@��#��@                        ��/���@H�4H�4@                H�4H�4@        ��/���@        ;��,��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#��@                        ��/����?0#0# @        ��/����?                        0#0# @;��,��@��/����?                ��/����?        ;��,��@                ;��,��@        0#0# @��#���?        0#0# @��#���?                                0#0# @��#��@                ��b:��*@��/����?H�4H�4@;��,��$@��/����?H�4H�4@;��,��$@��/����?0#0#�?��#�� @��/����?0#0#�?��#�� @��/����?                ��/����?        ��#�� @��/����?                ��/����?        ��#�� @                                0#0#�?��#�� @                ��#�� @                z�5��@                                0#0# @z�5��@                Mp�}N@t�'�x�R@5#0#`@��b:��:@��On�H@]��Y��X@��b:��:@��h
�G@��)��)C@<��,��4@��]�ڕE@��-��-5@        ��/���>@�C=�C=,@        Nn��O0@H�4H�4(@        0����/#@0#0#�?        �cp>@                ��/���@0#0#�?                0#0#�?        ��/���@                ���-��@#0#0&@        ���-��@0#0#@        ��/���@0#0#@        ��/���@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        �cp>@                        H�4H�4@        �cp>@                        �C=�C=@        ��|��,@0#0# @                0#0# @        ��|��,@        <��,��4@��On�(@�C=�C=@��#�� @/����/#@                D�JԮD!@                ��/����?                ���-��@        ��#�� @��/����?        ��#�� @                        ��/����?        �k(��2@�cp>@�C=�C=@�P^Cy/@        0#0#�?��#���?        0#0#�?��#���?                                0#0#�?���>��,@                z�5��@�cp>@H�4H�4@z�5��@                        �cp>@H�4H�4@        ��/����?H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@                H�4H�4@        ��/����?        z�5��@��/���@S2%S2%1@z�5��@��/���@S2%S2%1@z�5��@�cp>@0#0# @        �cp>@0#0#�?        ��/����?                ��/����?0#0#�?                0#0#�?        ��/����?        z�5��@        0#0#�?                0#0#�?z�5��@                        ��/����?�A�A.@        ��/����?H�4H�4@                H�4H�4@        ��/����?                        vb'vb'"@z�5��@                        �cp>@�A�AN@                �
��
�E@        �cp>@S2%S2%1@        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?0#0#0@                �A�A.@        ��/����?0#0#�?        ��/����?                        0#0#�?��#��@@�cp>�9@�A�A>@��#���?鰑%@0#0# @��#���?E�JԮD!@H�4H�4@                H�4H�4@��#���?D�JԮD!@        ��#���?��/����?                ��/����?        ��#���?                        ���-��@                ��/����?��+��+@        ��/����?                        ��+��+@���b:@@��/���.@#0#06@���b:@@���-��*@��+��+@���b:@@鰑%@��+��+@+�����;@0����/@��+��+@,�����;@��/����?��+��+@��#��@��/����?H�4H�4@        ��/����?        ��#��@        H�4H�4@z�5��@                ��#���?        H�4H�4@��#���?        0#0#�?                0#0#�?��#���?                                0#0# @�,����7@��/����?0#0# @        ��/����?        �,����7@        0#0# @������3@                ��#��@        0#0# @                0#0# @��#��@                        �cp>@                ��/����?                ��/����?        ��#��@�cp>@        z�5��@��/����?                ��/����?        z�5��@                ��#���?0����/@        ��#���?                        0����/@                �cp>@                ��/����?                ��/����?                ��/����?S2%S2%1@                ��+��+$@        ��/����?�C=�C=@                H�4H�4@        ��/����?0#0#@        ��/����?0#0#�?        ��/����?                ��/����?0#0#�?                0#0#�?        ��/����?                        H�4H�4@��#�� @��/����?0#0#0@��#�� @        H�4H�4@                0#0# @��#�� @        0#0#�?��#�� @                                0#0#�?        ��/����?��8��8*@        ��/����?                        ��8��8*@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ1�.hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKŅ�h��B+         l                 @�A�?��vbH�?#      M�t}@       [                 �|F�?*�����?�       _�\ؿj@                         ����?����L�?|       ��g��g@                        �q�3?0D>��?       �x4E@                           �?
4=�%�?       6���8@                        ,*�����?       ��l}�'*@                        �5W�?��|��?       ���ĺw@                        �YV?
4=�%�?       �(J��@	       
                 �dW?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               ��/����?������������������������       �      м       ��/����?������������������������       �               z�5��@                         
?�@ȱ��?	       nm���S'@                       ���I?�^�#΀�?       O�{��A%@������������������������       �               ��#���?                        ���i?      �<       0����/#@������������������������       �               ��/����?������������������������       �               ��/���@������������������������       �      �<       ��#���?                        fR�8?      �<       E�JԮD1@������������������������       �               ��/���@������������������������       �        
       ���-��*@       Z                 @4�?j������?]       l%H���b@       =                 PeT�?L2�$[�?Y       � Qt�a@       :                 p�x�?�̨r�{�?;       ��-<�V@       7                 ���?�~��.��?5       �EJ�T@       .                  �~��?�����?,       }$S��Q@       +                 ���z?:<��?       *:M_Z�4@       &                  �P��?,�^��?       A<��*�2@        #                 @F��3���r�?
       ��7�nN*@!       "                 P� ?� �_rK�?       J�@��"@������������������������       �               ;��,��@������������������������       �      ��       ��/���@$       %                 �p}?      �<       ��#��@������������������������       �               ��#���?������������������������       �               z�5��@'       (                  �a�?|@ȱ��?       nm���S@������������������������       �      ��       ��/���@)       *                   s��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?,       -                 �6�?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?/       6                 �y���@��K��?       ���0�H@0       3                 �T?�x�<�?
       X&b��q1@1       2                   �x�?ܗZ�	7�?       i~���@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?4       5                 �B{s?      �<       z�5��(@������������������������       �               z�5��@������������������������       �               �k(��"@������������������������       �               ���b:@@8       9                 �"c?,%@�"�?	       ��[�'@������������������������       �               ��/���@������������������������       �               ��#��@;       <                 p�f�?�5JH���?       �MOI#@������������������������       �               E�JԮD!@������������������������       �               0#0#�?>       W                 �ۙ�?_���1�?       e�&v�H@?       P                 ��{�? �ѩ<�?       &	��SB@@       E                  P�"�?��z}-�?       ��(�I�9@A       B                  [U�?�ۜ�x�?       d��إV#@������������������������       �      ȼ       ���-��@C       D                 �Iݩ?h%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?F       O                 ����?h�p����?       T�Ĭ�G0@G       N                 ���?�B���?       F��,�,@H       M                 �.��?
4=�%�?       �(J��@I       J                 0vb�?Ȕfm���?       ��Z�N@������������������������       �               ��#���?K       L                  `���?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ȼ       �k(��"@������������������������       �               0#0# @Q       V                 k�!?Z�ђ���?       �oFݜh%@R       U                    �? 4=�%�?       �(J��@S       T                  '�?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               �cp>@X       Y                 �R�־�o����?       ���5u*@������������������������       �               �cp>@������������������������       �      �<       <��,��$@������������������������       �               ���>��@\       c                 @5�?���?       F�X�U�6@]       `                 ����?���A���?       ��\�F"@^       _                 P��;?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?a       b                 �6�?��ڰ�x�?       �K�f�@������������������������       �               ;��,��@������������������������       �               0#0#�?d       e                 H{e�?�Qk��?       ��Th!�+@������������������������       �               0#0#@f       k                  �g<�?h�4���?       �tCP��#@g       j                    �?�;�a
=�?       ��l��@h       i                  X��?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?������������������������       �               ��/���@������������������������       �               H�4H�4@m       �                 @��?��T֙�?�       gɳ�2p@n       �                 ���c?@��#7��?       :��xuC@o       x                 ���s?*cL��?       ��Y|p�=@p       q                  ��?dV�\Ga�?
       q�6t%@������������������������       �               0#0#�?r       s                 �$��?b%��̫�?	       �@�o#@������������������������       �               ��/���@t       u                 ��x�?��íxq�?       $2��-�@������������������������       �      ��       ��/���@v       w                 �\2�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?y       �                 ԰�C?𜋙��?       aJ9U63@z                        �Q�?�d�$���?	       <��#�.@{       ~                 ��~?����X��?       &��֞&@|       }                ���c?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       �k(��"@�       �                 P���?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @�       �                 aؑ?̔fm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@�       �                 ܇�?x����?       �����!@������������������������       �               ��+��+@�       �                 Pl?x�G���?       ��%�|@������������������������       �               0#0#�?�       �                  2�i?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                  �g<�?�:��B�?~       �d�Kk@�       �                  �9��?g��|?�?!       �,��>J@�       �                 mm?�m��u;�?       ��5t@@�       �                 ����?�[�?$�?       :ha��7@�       �                 �yFC?���;�1�?       �$�S՞1@�       �                 ��?��
+���?	       \Zz�+�#@�       �                 �e_�?�26�
�?       4��*8E@�       �                 ���?�djH�E�?       ^�\m�n@�       �                 �I}�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?�       �                    �?����?       ��X�)B@������������������������       �               ��#�� @�       �                 `s5�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ȼ       ��/����?������������������������       �      Լ       �cp>@������������������������       �      ��       ��/���@������������������������       �      ȼ       z�5��@������������������������       �               vb'vb'"@�       �                 �zb�?`�4���?
       �tCP��3@������������������������       �               �cp>'@������������������������       �               0#0# @�       �                   ��?6֨�wO�?]       ��{e�d@�       �                 ����?�]?�?3       0%x�_U@�       �                 (�to?p�0���?       ���ϝ@@�       �                   �x�?a$�*��?       M{���2@�       �                    �?�/KI$��?       B��t&@������������������������       �               z�5��@�       �                   (�?f,���O�?       ���/> @������������������������       �               H�4H�4@������������������������       �               ��#�� @������������������������       �      �<       ��/���@������������������������       �               ��8��8*@�       �                 �O�?p���o�?       �SXOa�J@������������������������       �               ~˷|˷I@�       �                  `�J�?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?�       �                 �|'�?b��`p��?*       Ӣ9hKT@�       �                 �DF�?���!��?       sCP��H@������������������������       �               0����/@�       �                  ~�?x�G���?       ��ɘ�E@�       �                  �Ԧ�?��[����?       Gl�_A;@�       �                 �H��?���d��?       ��GQ�-@�       �                  �~��?���};��?       ��;̑�%@������������������������       �               �cp>@������������������������       �               0#0# @������������������������       �      �<       ��/���@������������������������       �               ��On�(@�       �                 @8��?w�;B��?	       ՟���	0@������������������������       �               H�4H�4(@�       �                 �$I�?x�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               0#0#@@�t�bh�hhK ��h��R�(KK�KK��h �Bx  ��tӹa@�����d@�ڬ�ڬd@
��G�[@I��t��V@H�4H�4(@2����"Z@^�ڕ��T@H�4H�4@<��,��$@�]�ڕ�?@        ;��,��$@��|��,@        ��#�� @0����/@        ��#�� @0����/@        ��#�� @�cp>@        ��#�� @��/����?                ��/����?        ��#�� @                        ��/����?                ��/����?        z�5��@                ��#�� @0����/#@        ��#���?/����/#@        ��#���?                        0����/#@                ��/����?                ��/���@        ��#���?                        E�JԮD1@                ��/���@                ���-��*@        �t�Y�W@�cp>�I@H�4H�4@�k(���U@�cp>�I@H�4H�4@�P^CyO@��|��<@0#0#�?�P^CyO@&jW�v%4@        ���>��L@��On�(@        ;��,��$@鰑%@        <��,��$@E�JԮD!@        �k(��"@��/���@        ;��,��@��/���@        ;��,��@                        ��/���@        ��#��@                ��#���?                z�5��@                ��#���?0����/@                ��/���@        ��#���?��/����?        ��#���?                        ��/����?                ��/����?                ��/����?                ��/����?        �,����G@��/����?        �P^Cy/@��/����?        z�5��@��/����?        z�5��@                        ��/����?        z�5��(@                z�5��@                �k(��"@                ���b:@@                ��#��@��/���@                ��/���@        ��#��@                        D�JԮD!@0#0#�?        E�JԮD!@                        0#0#�?|�5��8@�cp>7@0#0# @���>��,@&jW�v%4@0#0# @z�5��(@�cp>'@0#0# @��#���?E�JԮD!@                ���-��@        ��#���?��/����?        ��#���?                        ��/����?        \Lg1��&@�cp>@0#0# @[Lg1��&@�cp>@        ��#�� @�cp>@        ��#���?�cp>@        ��#���?                        �cp>@                ��/����?                ��/����?        ��#���?                �k(��"@                                0#0# @��#�� @E�JԮD!@        ��#�� @�cp>@        ��#���?�cp>@        ��#���?                        �cp>@        ��#���?                        �cp>@        ;��,��$@�cp>@                �cp>@        <��,��$@                ���>��@                z�5��@��/���@vb'vb'"@z�5��@��/����?0#0#�?��#���?��/����?                ��/����?        ��#���?                ;��,��@        0#0#�?;��,��@                                0#0#�?        �cp>@0#0# @                0#0#@        �cp>@0#0#@        �cp>@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/���@                        H�4H�4@�P^Cy?@>l��F:R@��)��)c@���>��,@��/���.@vb'vb'"@���>��,@���-��*@0#0# @��#���?��/���@0#0# @                0#0#�?��#���?��/���@0#0#�?        ��/���@        ��#���?��/���@0#0#�?        ��/���@        ��#���?        0#0#�?��#���?                                0#0#�?��b:��*@�cp>@        z�5��(@�cp>@        <��,��$@��/����?        ��#���?��/����?                ��/����?        ��#���?                �k(��"@                ��#�� @��/����?                ��/����?        ��#�� @                ��#���?�cp>@        ��#���?                        �cp>@                ��/����?�C=�C=@                ��+��+@        ��/����?0#0# @                0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?        ��#��0@��|��L@u�qb@<��,��$@�e�_��7@vb'vb'2@<��,��$@��On�(@��+��+$@;��,��$@��On�(@0#0#�?��#��@��On�(@0#0#�?��#��@0����/@0#0#�?��#��@��/����?0#0#�?��#��@��/����?0#0#�?��#���?        0#0#�?��#���?                                0#0#�?z�5��@��/����?        ��#�� @                ��#���?��/����?        ��#���?                        ��/����?                ��/����?                �cp>@                ��/���@        z�5��@                                vb'vb'"@        �cp>'@0#0# @        �cp>'@                        0#0# @z�5��@�-����@@I`F`�_@z�5��@��/���@n�fm��Q@;��,��@��/���@��)��)3@;��,��@��/���@H�4H�4@;��,��@        H�4H�4@z�5��@                ��#�� @        H�4H�4@                H�4H�4@��#�� @                        ��/���@                        ��8��8*@��#���?        ��8��8J@                ~˷|˷I@��#���?        0#0#�?                0#0#�?��#���?                        �cp>�9@�;�;K@        �cp>�9@#0#06@        0����/@                鰑5@#0#06@        /����/3@0#0# @        ���-��@0#0# @        �cp>@0#0# @        �cp>@                        0#0# @        ��/���@                ��On�(@                ��/����?�C=�C=,@                H�4H�4(@        ��/����?0#0# @        ��/����?                        0#0# @                0#0#@@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJg�)hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKh��BH4         �                 ��?���XT�?(      �)_a�}@       �                  �h?�'!h	s�?�       ˤgD�s@       �                 ��H?�	�{�?�       �A�m
Ip@       {                  `<��?���o�?�       8Λ糫k@       r                 ��@�?w<��,��?       h�y�i@       q                  `��?�)�[��?u       �6(���f@       Z                   �0�?r0���?p       V���e@       1                  �P��?��I��?`       ݕ� /�b@	       0                 �C>?��X���?.       �s����R@
                        ���>�l��?*       -5��tsQ@������������������������       �               ;��,��@                        �5�	?z�&�m��?'       x��:(P@                        @.��>Ȕfm���?       ��Z�N@                         
?\n����?       � ��w<@                        �؉�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#���?������������������������       �               0����/@       +                 ���?lG�m��?"       �ۉ��fL@                         ��^�?~�����?       ���/�D@������������������������       �               ��/����?                        �b�c?v���S~�?       �{��C@                        �#h?�N:�*ط?
       I�G�3@������������������������       �        	       �k(��2@������������������������       �      �<       ��/����?                        �O��?(mQ����?       ��1��K4@������������������������       �               ��/����?                         �u��?d���q�?       ��~�`2@������������������������       �               ��/����?                          o[?Х��Y��?       �u%!!k1@������������������������       �               ��/����?!       &                   ҏ�?��s`���?
       ���1�u0@"       %                    �?����?       ��X�)B@#       $                 �)88?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               ��#���?'       *                 �[�Z?��+%�"�?       ��kw��(@(       )                 h�&r?L� P?)�?       ����x�@������������������������       �               0#0#�?������������������������       �               ��#��@������������������������       �               ���>��@,       /                 �q�3?R��h���?       k��:�-@-       .                 ��}�?���Ѯ�?       ��GQ&@������������������������       �               �cp>@������������������������       �               ��#�� @������������������������       �      ȼ       ��/���@������������������������       �      �       �cp>@2       Q                 �(+�?��v��?2        �G.��R@3       B                 pb!i?0-Hg��?'       fo�+EM@4       ?                 �7�<?�7�֥��?       0����-?@5       >                 PGT~?���/��?       @z$S��7@6       =                    �?
4=�%�?       �(J��3@7       <                 �1�?�)z� ��?
       �\�,@8       ;                 �0��>�d�$���?       �T�f$@9       :                 p���?���/��?       V��7�@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      �<       z�5��@������������������������       �      ȼ       ��/���@������������������������       �      ��       �cp>@������������������������       �               ��#��@@       A                 ���A?      �<       ���>��@������������������������       �               ��#���?������������������������       �               z�5��@C       J                 p�%h?��n��?       �-H�\;@D       I                 �uY�?������?       �0G��l2@E       F                 ?}|?����VV�?	       A�R.�.@������������������������       �               ��On�(@G       H                 �m�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               H�4H�4@K       L                 �S�t?>�c3���?       �uk��!@������������������������       �               z�5��@M       N                  Ц6�?r@ȱ��?       om���S@������������������������       �               ��/���@O       P                 ��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?R       Y                 �;��?ߝ  ~�?       P@��W1@S       T                 \�ԑ?DF�X��?
       .�=k�U0@������������������������       �               z�5��@U       X                 ���?hP�D�?       �A��P?$@V       W                 �2*�?F���'0�?       �C�� T"@������������������������       �               ��/����?������������������������       �      ��       ���>��@������������������������       �      м       ��/����?������������������������       �               0#0#�?[       j                  `%+�?���(��?       B.�0~6@\       g                    �?8ĩAf�?       ��d>v�0@]       f                 X��3?hSmd�d�?       :��P{�@^       e                 ���?��r�g��?       ��1ֻ�@_       d                 �{�?����]L�?       N66�ͯ@`       c                 ���p?Ȕfm���?       ��Z�N@a       b                   ���?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �      м       ��/����?h       i                 �?      �<       D�JԮD!@������������������������       �               �cp>@������������������������       �               �cp>@k       l                 h'v�?���/��?       @z$S��@������������������������       �               ��#�� @m       n                 �۶�?Ȕfm���?       ��Z�N@������������������������       �               ��/����?o       p                 x!j�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#�� @s       z                  ���?x+}1�?
       �Vc��2@t       y                 p���?x��y�a�?	       +��lL/@u       v                 ��_�?����*�?       �	�c/(+@������������������������       �               ���-��@w       x                 �q��?�w��d��?       �0���s@������������������������       �               ��/���@������������������������       �      �<       H�4H�4@������������������������       �               ��#�� @������������������������       �               H�4H�4@|       �                 `#��?�3��F��?       nf9t{y4@}       �                 8݀t?$#����?       x�߄�3@~                        `$�a?`n����?       � ��w<@������������������������       �               ��#��@������������������������       �      �<       ��/����?�       �                 ؘl�?      �<       ��b:��*@������������������������       �               ��#�� @������������������������       �               ZLg1��&@������������������������       �      �<       ��/����?�       �                 `�??�����+�?       V�Ѓ�C@�       �                 ����?��q�R�?       �]�{�"@�       �                 �|L?z�G���?       '5L�`�@������������������������       �               ��/����?�       �                 �Ԇ�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               z�5��@�       �                 ����?���L
��?       ��e�0>@�       �                 0�Y? � N��?       �L�EBC3@������������������������       �               ��#���?������������������������       �               :l��F:2@�       �                  Ц6�?V����?       �Y9��%@������������������������       �               0����/@�       �                 ̤�?�J���?       a���@������������������������       �               z�5��@������������������������       �               H�4H�4@�       �                 �8U|?�τ%&�?       >��>F@�       �                 '�Ki?z��`p��?       �����@������������������������       �               ��/����?������������������������       �      ��       0#0#@�       �                 x�׀? �ދ��?       :UF#C@�       �                 P�J�?v=���?       � ��R(@������������������������       �               ��/����?������������������������       �               #0#0&@������������������������       �      ��       ��8��8:@�       �                  t�?h7����?g       g
�9��d@�       �                 �E�e?��ɰ��?E       �i�B]@�       �                 0�,�?`���
��?-       �?��/nR@������������������������       �               ;��,��$@�       �                 �jU?t�"J:�?'       �pv�O@�       �                 @�r�?&�Hx��?$       c�H��SL@������������������������       �               ��/���@�       �                ��G�?�=C:5�?"       u�˲hJ@�       �                 <�Q?T�n���?       K�D�I:@�       �                  ;��?��)|���?       ��R^7@�       �                 ���?�����?       �}WU0�2@�       �                    �?R��]H��?       ��v 1@�       �                 �rT�?8 d�?       "�ѿ-$@������������������������       �               ��+��+@�       �                 0��?ҟ��X�?       l�n�/@������������������������       �               0#0# @�       �                 ����?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?�       �                 @�#�?�AP�9��?       i��6��@������������������������       �               0#0#@�       �                  �3��?�� ��?       rp� k@������������������������       �               ��/����?�       �                 �zN�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      м       ��/����?�       �                 �j%?      �<       ��#��@������������������������       �               ��#�� @������������������������       �               ��#�� @�       �                 �^7�?b%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 `s5�?�L�ú��?       �����:@�       �                  н��?�Qk��?       ��Th!�@������������������������       �               �cp>@������������������������       �               0#0#@�       �                  `��?� {v�J�?       /��}��3@�       �                 p
E�?����?       ���"�X$@�       �                 ���?��t1u�?       "�te!� @�       �                 X�:�?�zœ���?       IG���t@������������������������       �               z�5��@������������������������       �               0#0#�?������������������������       �      ��       ��#��@������������������������       �      ȼ       ��/����?�       �                 @C��?ܜ�x�?       d��إV#@������������������������       �               ��/���@�       �                 �ec�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                  ��?      �<       ���-��@������������������������       �               ��/���@������������������������       �               �cp>@�       �                 �Ys�? ~�; -�?       Z��־�E@������������������������       �      м       0#0#@@�       �                 �C+�?�^�F�M�?       ��ޚ�&@������������������������       �               ��+��+$@������������������������       �      ȼ       ��/����?�       �                 Б0�?�Z� 5�?"       ���jI@�       �                  ���?�m��.�?        �xK&�H@������������������������       �               �cp>@�       �                  ��?� 	�?       T:E?n�F@�       �                  y��?|��`p��?       �����@������������������������       �               0#0# @�       �                 �'�?|�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 �@�?�2t �?       [�	v�C@������������������������       �               �s?�s?=@�       �                 �C8�?�o���?       p�9�F$@������������������������       �               ��#���?�       �                 ��^?l���X��?       Pà4�4"@�       �                 ،��?�o���?       o�9�F@������������������������       �               ��#���?������������������������       �               0#0#@�       �                8w}f�?      �<       0#0#@������������������������       �               0#0#�?������������������������       �               H�4H�4@�       �                 �h��?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?�t�bh�hhK ��h��R�(KK�KK��h �Bh  y�YLGc@�z����c@��+��+d@'�}��_@�����]@�A�AN@&�}��_@��|��\@��)��)3@+���>�]@���|NV@��8��8*@�}�\Y@��]�ڕU@��8��8*@�5��X@s�'�x�R@�C=�C=@^Lg1��V@r�'�x�R@�C=�C=@����bzU@�_��e�M@H�4H�4@6��tSH@�cp>�9@0#0#�?4��tSH@%jW�v%4@0#0#�?;��,��@                �k(���E@(jW�v%4@0#0#�?��#�� @�cp>@        ��#�� @��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#���?                        0����/@        =��,��D@��|��,@0#0#�?��#��@@��/���@0#0#�?        ��/����?        ��#��@@�cp>@0#0#�?�k(��2@��/����?        �k(��2@                        ��/����?        ���>��,@0����/@0#0#�?        ��/����?        ���>��,@�cp>@0#0#�?        ��/����?        ���>��,@��/����?0#0#�?        ��/����?        ���>��,@��/����?0#0#�?z�5��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ��#���?                [Lg1��&@        0#0#�?��#��@        0#0#�?                0#0#�?��#��@                ���>��@                ��#�� @���-��@        ��#�� @�cp>@                �cp>@        ��#�� @                        ��/���@                �cp>@        �k(��B@�-����@@��+��+@�,����7@��/���>@0#0#@������3@�cp>'@        z�5��(@�cp>'@        ��#�� @�cp>'@        ��#�� @�cp>@        ��#�� @��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        z�5��@                        ��/���@                �cp>@        ��#��@                ���>��@                ��#���?                z�5��@                ��#��@0����/3@0#0#@        ��|��,@0#0#@        ��|��,@0#0#�?        ��On�(@                ��/����?0#0#�?                0#0#�?        ��/����?                        H�4H�4@��#��@0����/@        z�5��@                ��#���?0����/@                ��/���@        ��#���?��/����?        ��#���?                        ��/����?        ��b:��*@�cp>@0#0#�?��b:��*@�cp>@        z�5��@                ���>��@�cp>@        ���>��@��/����?                ��/����?        ���>��@                        ��/����?                        0#0#�?;��,��@On��O0@0#0#�?��#�� @���-��*@0#0#�?��#�� @0����/@0#0#�?��#�� @�cp>@0#0#�?��#���?�cp>@0#0#�?��#���?�cp>@        ��#���?��/����?                ��/����?        ��#���?                        ��/����?                        0#0#�?��#���?                        ��/����?                D�JԮD!@                �cp>@                �cp>@        z�5��@�cp>@        ��#�� @                ��#���?�cp>@                ��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#�� @                ��#�� @鰑%@H�4H�4@��#�� @鰑%@H�4H�4@        鰑%@H�4H�4@        ���-��@                ��/���@H�4H�4@        ��/���@                        H�4H�4@��#�� @                                H�4H�4@��,���1@�cp>@        ��,���1@��/����?        ��#��@��/����?        ��#��@                        ��/����?        ��b:��*@                ��#�� @                ZLg1��&@                        ��/����?        ���>��@�cp>�9@H�4H�4@z�5��@�cp>@H�4H�4@        �cp>@H�4H�4@        ��/����?                ��/����?H�4H�4@        ��/����?                        H�4H�4@z�5��@                ��#��@�cp>7@H�4H�4@��#���?;l��F:2@        ��#���?                        :l��F:2@        z�5��@0����/@H�4H�4@        0����/@        z�5��@        H�4H�4@z�5��@                                H�4H�4@        �cp>@�ڬ�ڬD@        ��/����?0#0#@        ��/����?                        0#0#@        ��/����?�z��z�B@        ��/����?#0#0&@        ��/����?                        #0#0&@                ��8��8:@,�����;@2����/C@q�6k�6Y@�#���9@�]�ڕ�?@
����M@
�#���9@��/���>@S2%S2%1@;��,��$@                �P^Cy/@��/���>@S2%S2%1@�P^Cy/@�e�_��7@S2%S2%1@        ��/���@        �P^Cy/@%jW�v%4@S2%S2%1@���>��@���-��@H�4H�4(@z�5��@0����/@H�4H�4(@��#�� @0����/@H�4H�4(@��#�� @�cp>@H�4H�4(@��#�� @��/����?�C=�C=@                ��+��+@��#�� @��/����?0#0# @                0#0# @��#�� @��/����?        ��#�� @                        ��/����?                ��/����?��+��+@                0#0#@        ��/����?0#0#�?        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?        ��#��@                ��#�� @                ��#�� @                ��#���?��/����?        ��#���?                        ��/����?        ��#�� @���-��*@��+��+@        �cp>@0#0#@        �cp>@                        0#0#@��#�� @鰑%@0#0#�?���>��@��/����?0#0#�?���>��@        0#0#�?z�5��@        0#0#�?z�5��@                                0#0#�?��#��@                        ��/����?        ��#���?D�JԮD!@                ��/���@        ��#���?��/����?        ��#���?                        ��/����?                ���-��@                ��/���@                �cp>@                ��/����?��-��-E@                0#0#@@        ��/����?��+��+$@                ��+��+$@        ��/����?        ��#�� @���-��@�ڬ�ڬD@��#�� @0����/@�ڬ�ڬD@        �cp>@        ��#�� @��/����?�ڬ�ڬD@        ��/����?0#0#@                0#0# @        ��/����?0#0# @        ��/����?                        0#0# @��#�� @        �z��z�B@                �s?�s?=@��#�� @        0#0# @��#���?                ��#���?        0#0# @��#���?        0#0#@��#���?                                0#0#@                0#0#@                0#0#�?                H�4H�4@        ��/����?                ��/����?                ��/����?        �t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�]_AhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK���h��Bx(         �                 ��g?:�9��L�?      \O�k�w}@       u                 ��??���c��?�       �\�<�u@       n                 ���?�u���[�?�       ��L/5o@       W                 �^Ҧ?�>k�6��?�       �v�X�tl@       P                 ���?���.*!�?o       �剿�kg@       /                 �x�?�)�yt��?c       ^`Il��d@                        "?�뇑��?>       �Y�[@                        �y���HBms�?       ��֖��;@	       
                   �P�?��Z�	7�?       j~���@������������������������       �               ��#�� @                        ��?f%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?                        �Y֬>      �<       \Lg1��6@������������������������       �               ��#���?������������������������       �               �k(���5@                        P��i?��7m�?-       �(�+T@                        ��IL?fQ��?       �s�=�1@                        �3�_?�d�$���?       �T�f@                        ���?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               ��#�� @������������������������       �      ��       ��On�(@                        P�ϊ?J1`f+q�?"       6�W���O@                        �j[?P�F¯?       �:.�=@������������������������       �      ȼ
       ��,���1@                        ����?|b8�Y�?       FJͰ(@������������������������       �      �<       ZLg1��&@������������������������       �      ȼ       ��/����?       ,                 ����?�ԏj��?       �~:�.�@@        +                �3G�y?��w"T�?       �W����5@!       "                 `�ג?���'��?       �v�9��4@������������������������       �               D�JԮD!@#       *                 �j��?fn����?       � ��w<(@$       %                 ���j?X�j���?       ���z"@������������������������       �               ;��,��@&       )                    �?�����?       ��X�)B@'       (                 P#%v?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               ��#���?������������������������       �      ȼ       �cp>@������������������������       �               ��#���?-       .                  �.�?      �<       \Lg1��&@������������������������       �               ��#��@������������������������       �               ���>��@0       I                 ��^�?-����?%       pKr�� M@1       F                 P��?X�,��?       �t5ëF@2       E                      ^|*įS�?       q�go'@@3       @                    �?Fͻ�&��?       |���g�1@4       ?                  ����?���/��?	       @z$S��'@5       <                ��r?��Z�	7�?       j~���$@6       7                 �-�?���/��?       V��7�@������������������������       �               z�5��@8       ;                 `�p�?& k�Lj�?       �q��l}@9       :                 L�Q�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       �cp>@=       >                �va�?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?������������������������       �      ��       ��/����?A       B                  �]�?t@ȱ��?       om���S@������������������������       �               �cp>@C       D                ���c?b%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �      �<       ��|��,@G       H                 @���?�3���r�?       ��7�nN*@������������������������       �               ��/���@������������������������       �      ��       �k(��"@J       K                 P�s�?N0�8���?	       #Z��!�)@������������������������       �               �cp>@L       O                 ��B�?�?�0�!�?       a`�T�$@M       N                 GW�d?����|e�?       �z �B�@������������������������       �               H�4H�4@������������������������       �      �<       ��/����?������������������������       �               H�4H�4@Q       T                 `s��?0�#�Ѵ�?       �)�B�4@R       S                  �E�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @U       V                 X �?      �<
       ��,���1@������������������������       �               ��#���?������������������������       �        	       ��#��0@X       Y                 �V}?�lO��?       ^E�e�#D@������������������������       �               ��+��+@Z       i                 �I�?�S�g@�?       � V�A@[       h                 @8��?�f��m�?       ��OY>@\       g                 ���?��Oޤr�?       ��A�]=@]       b                  �Q�?
nw��?       b�?�-<@^       a                 p���?lSmd�d�?       :��P{�@_       `                 ��E�?T����1�?       ��;9�@������������������������       �               ��#�� @������������������������       �               0#0#�?������������������������       �               0����/@c       d                 �m�?�G�<�J�?       R �24@������������������������       �        	       ��|��,@e       f                 p���?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �               0����/@������������������������       �               0#0#�?������������������������       �      �<       ��#���?j       m                    �?�|2N��?       �3K}@k       l                 �5W�?�zœ���?       IG���t@������������������������       �               0#0#�?������������������������       �               z�5��@������������������������       �               0#0#�?o       p                  v�?.�O�:�?       �ʒ�6@������������������������       �               ��/����?q       t                 �_��?�IQ���?       ��]4@r       s                   �G�??�	,�?       >0�1b3@������������������������       �               ��/����?������������������������       �               S2%S2%1@������������������������       �      �<       ��#���?v       �                 ��+a?�
��?;       �\�*EX@w       �                 ���?8a_)��?!       e����J@x       �                 �P��?pC_}�O�?       ��0��D@y       ~                 ���?e��}�?       �|���BD@z       }                 ��vi?�4�A�?       �]j�,�A@{       |                 (I��?�^�#΀�?       P�{��A%@������������������������       �               /����/#@������������������������       �      �<       ��#���?������������������������       �               ��On�8@       �                 ��[�?4=�%�?       �(J��@������������������������       �               ��#�� @������������������������       �               �cp>@������������������������       �     ��<       0#0#�?�       �                 pM�D?�4��v�?	       �Y-"�'@������������������������       �               z�5��@�       �                 ��֬?lQ��?       �s�=�!@�       �                  ��G�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @�       �                    �?      �<       �cp>@������������������������       �               �cp>@������������������������       �               �cp>@�       �                 ���?-�؈��?       31��E@�       �                  `%+�?x�2|���?       �n�df_7@�       �                 е3g?�հ�.�?       �����X4@������������������������       �               ��#���?�       �                 �B��?�[nD���?       ���y�O3@�       �                 ��C?X%��̫�?       �@�o#@������������������������       �               0#0#�?�       �                  ~��?)���?       y��uk!@�       �                 ��0{?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ��       ���-��@������������������������       �               0����/#@������������������������       �               H�4H�4@�       �                  E(�?ֵ�d'�?       t����I4@�       �                 @��?����X��?       &��֞&@������������������������       �               �k(��"@�       �                 @� �?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 ���?l����?       �����!@������������������������       �               �C=�C=@������������������������       �      ȼ       ��/����?�       �                 �=�t?��+�c�?L       Rʫ�|/_@������������������������       �               ��#���?�       �                    �?�IuI�?K       .�=�^@������������������������       �        %       �C=�C=L@�       �                 @f�?�&��{�?&       <p���P@������������������������       �               �s?�s?=@�       �                 X�6�?j��e��?       z&[�}�B@�       �                 ����?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?�       �                 �C��?��i���?       ����A@������������������������       �               �A�A.@�       �                 ���o?��#���?       �͆�1�2@������������������������       �               H�4H�4@�       �                 Ј�v?B0�8���?	       "Z��!�)@������������������������       �               ��/����?�       �                  L��?��H�&p�?       L^�3��%@������������������������       �               ��/����?�       �                 �_��?�?�0�!�?       a`�T�$@������������������������       �               H�4H�4@�       �                 �Sl�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@�t�b�
     h�hhK ��h��R�(KK�KK��h �BX  �YLg1b@!jW�v%d@�ڬ�ڬd@�}��a@鰑Nc@H�4H�4H@���b:�^@�'�xr�V@vb'vb'B@��>���^@��]�ڕU@��)��)3@���>��\@2����-O@vb'vb'"@�5��X@��/���N@vb'vb'"@�b:���S@��|��<@        
�#���9@��/����?        z�5��@��/����?        ��#�� @                ��#���?��/����?                ��/����?        ��#���?                \Lg1��6@                ��#���?                �k(���5@                ��b:��J@���-��:@        ��#��@���-��*@        ��#��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ��#�� @                        ��On�(@        |�5��H@���-��*@        ���>��<@��/����?        ��,���1@                ZLg1��&@��/����?        ZLg1��&@                        ��/����?        <��,��4@��On�(@        �k(��"@��On�(@        ��#�� @��On�(@                D�JԮD!@        ��#�� @��/���@        ��#�� @��/����?        ;��,��@                z�5��@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ��#���?                        �cp>@        ��#���?                \Lg1��&@                ��#��@                ���>��@                ��#��0@Pn��O@@vb'vb'"@��#��0@��|��<@        ���>��@��On�8@        ���>��@鰑%@        z�5��@�cp>@        z�5��@��/���@        ��#��@��/���@        z�5��@                ��#���?��/���@        ��#���?��/����?                ��/����?        ��#���?                        �cp>@        ��#�� @                ��#���?                ��#���?                        ��/����?        ��#���?0����/@                �cp>@        ��#���?��/����?                ��/����?        ��#���?                        ��|��,@        �k(��"@��/���@                ��/���@        �k(��"@                        ��/���@vb'vb'"@        �cp>@                ��/����?vb'vb'"@        ��/����?H�4H�4@                H�4H�4@        ��/����?                        H�4H�4@������3@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ��,���1@                ��#���?                ��#��0@                z�5��@�e�_��7@��+��+$@                ��+��+@z�5��@�e�_��7@��+��+@z�5��@�e�_��7@H�4H�4@��#�� @�e�_��7@H�4H�4@��#�� @�e�_��7@0#0# @��#�� @0����/@0#0#�?��#�� @        0#0#�?��#�� @                                0#0#�?        0����/@                /����/3@0#0#�?        ��|��,@                0����/@0#0#�?                0#0#�?        0����/@                        0#0#�?��#���?                z�5��@        0#0# @z�5��@        0#0#�?                0#0#�?z�5��@                                0#0#�?��#���?��/���@S2%S2%1@        ��/����?        ��#���?��/����?S2%S2%1@        ��/����?S2%S2%1@        ��/����?                        S2%S2%1@��#���?                <��,��4@��P@H�4H�4(@��#�� @h
��F@0#0#�?z�5��@�+Q��B@0#0#�?z�5��@�+Q��B@        ��#���?F�JԮDA@        ��#���?0����/#@                /����/#@        ��#���?                        ��On�8@        ��#�� @�cp>@        ��#�� @                        �cp>@                        0#0#�?;��,��@���-��@        z�5��@                ��#�� @���-��@        ��#�� @��/����?                ��/����?        ��#�� @                        �cp>@                �cp>@                �cp>@        z�5��(@&jW�v%4@#0#0&@��#�� @D�JԮD1@0#0#@��#�� @E�JԮD1@0#0#�?��#���?                ��#���?E�JԮD1@0#0#�?��#���?��/���@0#0#�?                0#0#�?��#���?��/���@        ��#���?��/����?                ��/����?        ��#���?                        ���-��@                0����/#@                        H�4H�4@;��,��$@�cp>@�C=�C=@;��,��$@��/����?        �k(��"@                ��#���?��/����?                ��/����?        ��#���?                        ��/����?�C=�C=@                �C=�C=@        ��/����?        ��#���?���-��@�s?�s?]@��#���?                        ���-��@�s?�s?]@                �C=�C=L@        ���-��@�A�AN@                �s?�s?=@        ���-��@=�C=�C?@        �cp>@0#0#�?        �cp>@                        0#0#�?        ��/���@�A�A>@                �A�A.@        ��/���@�A�A.@                H�4H�4@        ��/���@vb'vb'"@        ��/����?                ��/����?vb'vb'"@        ��/����?                ��/����?vb'vb'"@                H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJL�OhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKم�h��Bx/         h                  �~��?N��V?@�?'      ��\��}@                        `�yS?�E`���?t       �;��|g@������������������������       �               鰑%@       I                 P7&E? �;k#�?n       ?-qf*f@                          �G�?��'qV��?M       �� `@                        �;�j?�z���`�?       �7���@@                         ��F&Μ�!�?	       D3�\r.@������������������������       �               ��/����?	       
                 0�3I?�(߫$��?       0H����*@������������������������       �               �k(��"@                        ���8?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @                        �Q�?B4|���?       �T|qt2@                        XFe�?�Tu��?       ����.@������������������������       �      �<       ��On�(@                         `�J�?^%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?                           �?hn����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?       F                 P�?�� U�?9       h�m�ٰW@       =                 pTF�?��~��?6       N,�5�V@       &                 ����?�H�o�?*       dy�DgR@                        ����?T�s�	�?       �rD@                        ~`���_�A�?       肵�e`@                        �NR?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               z�5��@        #                 ���a?0�#�ݬ?       0X{Z�@@!       "                 0�R�?�����?       �O��@������������������������       �               ;��,��@������������������������       �      ȼ       ��/����?$       %                 �ao�>      �<       ��b:��:@������������������������       �               ��#���?������������������������       �               
�#���9@'       0                    �?6f辭}�?       9꜊v�@@(       /                 A��?T��h���?
       j��:�-@)       .                 0���?\n����?	       � ��w<(@*       -                      j��H��?       v�I�@+       ,                 8^q�?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@������������������������       �               �cp>@������������������������       �      ��       ;��,��@������������������������       �      �<       �cp>@1       6                 P���?�qL�Ľ�?
       ;W�w�y2@2       5                 �/�?�Ʈ^���?       �.g���,@3       4                  �JV�?T����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �               ZLg1��&@7       :                   .p�?�3`���?       .�r��@8       9                 ,.l�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?;       <                 h��1?      �<       0#0# @������������������������       �               0#0#�?������������������������       �               0#0#�?>       ?                  h��?B��aB��?       ����2@������������������������       �               ��/���@@       E                  �g<�?"�b���?	       �GXvƒ,@A       D                 ����?��ڰ�x�?       �K�f�(@B       C                 @�C�?�J���?       ��*]Y@������������������������       �               ��#�� @������������������������       �               0#0# @������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?G       H                 �.�?     ��<       H�4H�4@������������������������       �               0#0#�?������������������������       �               0#0# @J       W                 �vs�?�~ ��?!       �P�%qH@K       V                 ���?��f^�|�?       ��S�^u@@L       O                    �?��K�m��?       S�D]�>@M       N                 �%N�?�G�<�J�?       S �24@������������������������       �               /����/3@������������������������       �               0#0#�?P       Q                 ���G?V�ђ���?       �oFݜh%@������������������������       �               ��#���?R       U                 ��{�?�ۜ�x�?       d��إV#@S       T                   s��?��fm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               0#0# @X       c                 P�9�?,��V�"�?       ��y���/@Y       \                 p��?�/y߃�?       ǁ\��((@Z       [                 ���?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?]       b                 �Q�?�N̸��?       �#�zY9$@^       _                 0�֪?�o���?       o�9�F@������������������������       �               0#0# @`       a                 Ш��?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?������������������������       �               ��+��+@d       g                 �c(�?�@G���?       hu��@e       f                 �?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               0#0#�?i       �                 pG�?l�����?�       ѭR���q@j       s                 �۾c?��Z�k�?6       �-�V�V@k       l                 �KdU?�q��/��?       h
��F@������������������������       �               �cp>@m       p                 ��Bh?�#�Ѵ�?       �)�B�D@n       o                 P�Ab?�_�A�?       肵�e`@������������������������       �      �<       ;��,��@������������������������       �      ȼ       ��/����?q       r                    �?      �<       Fy�5A@������������������������       �               ��b:��:@������������������������       �               ���>��@t       �                 �ܣ�?�F��4��?       	�%��F@u       �                    �?�5�G|��?       �z�g�lD@v       �                 P���?��Z�	7�?       ���`�$>@w       ~                 p�ŗ?�3���r�?       ��7�nN:@x       }                 ���?��k{��?	       `;�W� *@y       |                 `]j�?jP�D�?       �A��P?$@z       {                  ��?
4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @������������������������       �               ;��,��@������������������������       �      �<       �cp>@       �                 `�
E?�(߫$��?       2H����*@�       �                  `���?L���'0�?       �C�� T"@�       �                  �?Z%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               z�5��@������������������������       �               ��#��@�       �                 �N��?      �<       ��/���@������������������������       �               ��/����?������������������������       �               ��/����?�       �                 @�?�?f�ђ���?       �oFݜh%@�       �                 �:��?      �<       D�JԮD!@������������������������       �               ��/����?������������������������       �               ���-��@������������������������       �               ��#�� @�       �                 d��?      �<       ��+��+@������������������������       �               H�4H�4@������������������������       �               0#0# @�       �                 �HϽ?��+҉G�?}       �D�h8kh@�       �                 `��\?Flxe�?e       �|w��Gc@�       �                 �9��?��vid�?9       ?�œ[�T@�       �                 ���?Q;Iֵ�?        ����m�F@�       �                 0Q�x?�ŉZ�N�?       ����@@�       �                 �$܀?X#��3��?	       j��Ѝ�)@�       �                 �M��?������?       +�ǟf%@�       �                 �؉�?xLU���?       h�ҹ^�@������������������������       �               0#0#�?������������������������       �               ���-��@�       �                  'n�?z��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 @��u?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?�       �                 �j��?�� ��8�?       ¶h�|x4@�       �                 ԰�C?�3`���?       .�r��@�       �                �J��?�D#���?       �B�j@������������������������       �               0#0# @������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 ��ߢ?��s`���?       ���1�u0@������������������������       �      ��       |�5��(@�       �                  �Q�?r�T���?       ��e[�&@������������������������       �               ��#�� @�       �                 0?x�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 P��?<@�����?       \n\�/V)@������������������������       �               H�4H�4@�       �                 p�L�?x5JH���?       �MOI#@�       �                ��S��?�@G���?       hu��@������������������������       �               0#0#�?������������������������       �               �cp>@������������������������       �      ȼ       �cp>@�       �                 GW�d?>3[ ���?       �֗CIC@�       �                 �fQ?<��0���?       V��I�!;@������������������������       �               k�6k�69@������������������������       �      ȼ       ��/����?�       �                 �!�?n�/W�D�?	       ���z^�%@�       �                 @� ?�����?       �v�qp�!@�       �                  0Y��?�֪u�_�?       ��?�8@������������������������       �               0����/@������������������������       �               0#0#�?������������������������       �               H�4H�4@�       �                 �N��?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?�       �                 ��W�?�F�]v>�?,       �@)f�Q@�       �                 p��?@}/W�?)       ��8#�P@������������������������       �               ;�;�F@�       �                 �.K�?@L�0�h�?       l�e�3@�       �                 �=��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               S2%S2%1@�       �                 ��"�?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �               0����/@�       �                 ��~? �-Zc�?       ��L^�D@������������������������       �               �cp>@�       �                 ਮ�?HL�0�h�?       k�e�C@�       �                    �?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 �j��?Pʊs`�?       �	S\!B@�       �                 0�i�?v=���?       � ��R(@�       �                 ��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��+��+$@������������������������       �      ��       H�4H�48@�t�bh�hhK ��h��R�(KK�KK��h �BX  cCy��d@B�JԮDa@�fm�f�d@�#����U@�JԮDmS@#0#06@        鰑%@        �#����U@�-����P@#0#06@���#8U@����z�A@0#0# @���>��,@1����/3@        [Lg1��&@��/���@                ��/����?        [Lg1��&@��/����?        �k(��"@                ��#�� @��/����?                ��/����?        ��#�� @                z�5��@��/���.@        ��#���?��|��,@                ��On�(@        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ��,���Q@On��O0@0#0# @��,���Q@Nn��O0@��+��+@Lp�}N@鰑%@H�4H�4@�k(��B@�cp>@        ;��,��@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                z�5��@                ���b:@@��/����?        ;��,��@��/����?        ;��,��@                        ��/����?        ��b:��:@                ��#���?                
�#���9@                \Lg1��6@��/���@H�4H�4@��#�� @���-��@        ��#�� @��/���@        z�5��@��/���@        z�5��@��/����?                ��/����?        z�5��@                        �cp>@        ;��,��@                        �cp>@        ���>��,@��/����?H�4H�4@��b:��*@        0#0#�?��#�� @        0#0#�?                0#0#�?��#�� @                ZLg1��&@                ��#���?��/����?0#0# @��#���?��/����?        ��#���?                        ��/����?                        0#0# @                0#0#�?                0#0#�?;��,��$@�cp>@0#0# @        ��/���@        ;��,��$@��/����?0#0# @;��,��$@        0#0# @��#�� @        0#0# @��#�� @                                0#0# @��#�� @                        ��/����?                        H�4H�4@                0#0#�?                0#0# @z�5��@�]�ڕ�?@�C=�C=,@��#�� @�a#6�;@H�4H�4@��#�� @�a#6�;@0#0#�?        0����/3@0#0#�?        /����/3@                        0#0#�?��#�� @E�JԮD!@        ��#���?                ��#���?E�JԮD!@        ��#���?�cp>@                �cp>@        ��#���?                        �cp>@                        0#0# @��#���?��/���@#0#0&@��#���?��/����?��+��+$@        ��/����?0#0#�?        ��/����?                        0#0#�?��#���?        vb'vb'"@��#���?        0#0#@                0#0# @��#���?        0#0# @                0#0# @��#���?                                ��+��+@        �cp>@0#0#�?        �cp>@                ��/����?                ��/����?                        0#0#�?�b:���S@=��18N@vb'vb'b@Np�}N@��On�8@��+��+@������C@0����/@                �cp>@        ������C@��/����?        ;��,��@��/����?        ;��,��@                        ��/����?        Fy�5A@                ��b:��:@                ���>��@                <��,��4@&jW�v%4@��+��+@;��,��4@&jW�v%4@        �k(��2@�cp>'@        �k(��2@��/���@        ���>��@�cp>@        ���>��@�cp>@        ��#�� @�cp>@                �cp>@        ��#�� @                ;��,��@                        �cp>@        ZLg1��&@��/����?        ���>��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        z�5��@                ��#��@                        ��/���@                ��/����?                ��/����?        ��#�� @D�JԮD!@                D�JԮD!@                ��/����?                ���-��@        ��#�� @                                ��+��+@                H�4H�4@                0#0# @������3@����z�A@cF`�a@������3@��/���>@�Wx�W�Y@������3@��On�8@������C@��,���1@:l��F:2@��+��+$@��,���1@0����/#@H�4H�4@��#�� @��/���@H�4H�4@        ��/���@H�4H�4@        ���-��@0#0#�?                0#0#�?        ���-��@                ��/����?0#0# @        ��/����?                        0#0# @��#�� @                ��#���?                ��#���?                �P^Cy/@��/����?H�4H�4@��#���?��/����?0#0# @��#���?        0#0# @                0#0# @��#���?                        ��/����?        ���>��,@��/����?0#0#�?|�5��(@                ��#�� @��/����?0#0#�?��#�� @                        ��/����?0#0#�?        ��/����?                        0#0#�?        E�JԮD!@0#0#@                H�4H�4@        E�JԮD!@0#0#�?        �cp>@0#0#�?                0#0#�?        �cp>@                �cp>@        ��#�� @���-��@�s?�s?=@        ��/����?k�6k�69@                k�6k�69@        ��/����?        ��#�� @0����/@0#0#@        0����/@0#0#@        0����/@0#0#�?        0����/@                        0#0#�?                H�4H�4@��#�� @                ��#���?                ��#���?                        �cp>@2#0#P@        ��/����?Q��N��O@                ;�;�F@        ��/����?vb'vb'2@        ��/����?0#0#�?        ��/����?                        0#0#�?                S2%S2%1@        0����/@0#0#�?                0#0#�?        0����/@                0����/@vb'vb'B@        �cp>@                ��/����?wb'vb'B@        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?eJ�dJ�A@        ��/����?#0#0&@        ��/����?0#0#�?        ��/����?                        0#0#�?                ��+��+$@                H�4H�48@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ��lhFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK���h��B�(         �                 0�0�?�@z�P�?#      �D�[�}@       S                 `�ݍ?PZ3����?�       �����vt@       R                 `��?D������?�       c���
Ki@       A                 0G?�y��:{�?�       U��8�h@       0                 �U���2���?h       h=���:d@                         ��?>/ќ4>�?=       iG��*X@                         ͺO?:v�qb�?+       |�v�9SQ@                        �\͵?bdؗ��?       4d��8@	                          �x�?��k{��?	       `;�W� *@
                         h��?nP�D�?       �A��P?$@������������������������       �               ��/����?                        �@?F���'0�?       �C�� T"@                            �?      �<       ���>��@������������������������       �               ��#���?������������������������       �               z�5��@������������������������       �      �<       ��/����?������������������������       �      ȼ       �cp>@������������������������       �               �cp>'@                        �
o?������?       [d�R�dF@                        �vs?���5�?       E�)�B=@                        ��h?�C=+��?
       b��T|0@������������������������       �               {�5��(@                         Џ~�?����?       ��X�)B@������������������������       �      ��       z�5��@������������������������       �      �<       ��/����?                        �C8�?0µ*A
�?
       ��A抌)@������������������������       �               ��#��@������������������������       �      ��       D�JԮD!@������������������������       �               �P^Cy/@       '                    �?:���@�?       �CA�9[;@       "                 ��H�?��$�|x�?       z"K�_:0@        !                h�ȼZ?b,���O�?       ���/>@������������������������       �               ��#���?������������������������       �               H�4H�4@#       $                  �_�?֬ͅV�?	       c�U(@������������������������       �               �cp>@%       &                 �W��?�wV����?       Bi�i�"@������������������������       �               ��#�� @������������������������       �               0#0#�?(       )                   E(�?E��I��?       �B��A&@������������������������       �               0#0#@*       /                 ���~?�_�A�?       炵�e`@+       .                 ��~?�����?       �O��@,       -                   ��?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               z�5��@������������������������       �      ȼ       ��/����?1       :                 �堘?�mÔx��?+       c3ˡ�KP@2       9                  ����?&�b�H�?$       ��~:��K@3       4                  y��?Zn����?       ����45@������������������������       �      ؼ	       ZLg1��&@5       8                 � 5?������?       �4^$4�#@6       7                 0��"?�����?       ��X�)B@������������������������       �               ��/����?������������������������       �      �<       z�5��@������������������������       �      ȼ       �cp>@������������������������       �               Ey�5A@;       <                 H�q?������?       �4^$4�#@������������������������       �               ��#�� @=       >                 `�m�?p�r{��?       e�6� @������������������������       �               ��/���@?       @                 p��?Ɣfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?B       Q                 @���?�sP�M=�?       ��H�B@C       L                  `���?�`���?       �f��/A@D       K                  gm?�j �N�?       y��4^6@E       J                 �.�\?�3+�Pr�?       Y-"�=L4@F       I                    �?Ȕfm���?       ��Z�N@G       H                 Pq8�?d%@�"�?       ��[�@������������������������       �      �<       ��/���@������������������������       �               ��#�� @������������������������       �               ��/����?������������������������       �      �<       ��On�(@������������������������       �      ܼ       ��#�� @M       N                 p'�H?Ny��]0�?       ���y"(@������������������������       �               ��/����?O       P                 �Q�?�^�F�M�?       ��ޚ�&@������������������������       �               ��/����?������������������������       �               ��+��+$@������������������������       �      �<       z�5��@������������������������       �      �       H�4H�4@T       a                  �g<�?�4��.�?K       �3�R�E_@U       \                 �U��>�Q��Ab�?       o��;@@V       [                  18�?�_�A�?
       悵�e`,@W       Z                  �?� �_rK�?       J�@��"@X       Y                 p���?�����?       �O��@������������������������       �               ��/����?������������������������       �      �<       ;��,��@������������������������       �               �cp>@������������������������       �               ;��,��@]       ^                 �8D�?�-����?       hM��F2@������������������������       �        
       ��/���.@_       `                   �G�?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?b       �                 ����?J�!Id�?5       �;�(W@c       |                 ��"}?�������?/       �7�bT@d       y                 p�7[?�1Qn�/�?%       6z��u�O@e       v                 GW�d?�y2cs�?       �����G@f       s                 ����?2rG�P��?       <|v-�D@g       r                 ���?�j��?       ��1g�4@h       q                  �E�?�!A_!�?       E����0@i       p                 B{�?�
�CX�?       ��:.�%@j       m                 ����?�y��d��?       �=�0�@k       l                  .s�?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@n       o                 @�w�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ��       ��/���@������������������������       �      ��       �cp>@������������������������       �               0#0#@t       u                 �\͵?      �<       ��-��-5@������������������������       �               0#0# @������������������������       �               ��)��)3@w       x                 �ңu?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/���@z       {                 �-�?      �<       0#0#0@������������������������       �               H�4H�4@������������������������       �               ��8��8*@}       �                 PFe�?���ج1�?
       ��+"6�1@~       �                 pO�v?灸�V/�?       ����|
*@       �                    �?���/��?       V��7�@������������������������       �               ��#��@������������������������       �      �<       ��/���@������������������������       �               ��+��+@������������������������       �               0����/@�       �                  P�"�?      �<       #0#0&@������������������������       �               0#0# @������������������������       �               vb'vb'"@�       �                 pJ�q?�>i��?W       S2���"b@�       �                 0�?��K�#�?+       g4N�%5Q@������������������������       �               ��b:��*@�       �                 ��C?������?'       (�h�K@�       �                 @� ?��5���?       �6��|A@�       �                 �I��?&��5�?       ��~���5@�       �                 H�6�?fm���?       �0��z'@�       �                 ��5�?R�ђ���?       �oFݜh%@������������������������       �               ��#�� @������������������������       �      ��       D�JԮD!@������������������������       �      ܼ       ��#���?�       �                 �W�?�i^�c�?       �D9�V$@������������������������       �               ;��,��@�       �                 4w�?�@����?       ���a�@�       �                 ����?z��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?������������������������       �               0#0# @�       �                 �;��?���<�?       f�W�l(@�       �                 0*tC?�~�Hs=�?       ��?Z[ @�       �                 tم�?\����?       P	K��@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?������������������������       �               0#0#�?������������������������       �               0#0#@�       �                 �`��?����A�?       ���,�@5@�       �                 ���? ����o�?       ^���v<3@������������������������       �        	       ��/���.@�       �                 Pj��?�@G���?       hu��@������������������������       �               0#0#�?�       �                 `�/S?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               0#0# @�       �                 �|'�??�	,�?,       >0�1bS@�       �                 �p�?�C��O�?       4�V��@@�       �                 P��?���L�?       >G���@@�       �                  �i�?D0�8���?       #Z��!�)@�       �                 ��=�?�w��d��?       �0���s@������������������������       �      �<       H�4H�4@������������������������       �               ��/���@������������������������       �               H�4H�4@�       �                 `�4x?L�0�h�?	       k�e�3@�       �                  0p��?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �      ��       0#0#0@������������������������       �      �<       ��/����?�       �                 ����?�n	�/��?       H�YŦ'E@������������������������       �      м       �A�A>@�       �                 ��ӣ?Dv=���?       � ��R(@������������������������       �               ��/����?������������������������       �               #0#0&@�t�bh�hhK ��h��R�(KK�KK��h �B�  �>��d@��e�_�b@�N��Nld@��#��`@����\@�ڬ�ڬT@���>��\@Rn��OP@��-��-5@���>��\@Rn��OP@vb'vb'2@��+[@�'�xr�F@0#0# @u�}wL@�]�ڕ�?@0#0# @���#8E@���-��:@        ���>��@D�JԮD1@        ���>��@�cp>@        ���>��@�cp>@                ��/����?        ���>��@��/����?        ���>��@                ��#���?                z�5��@                        ��/����?                �cp>@                �cp>'@        ��,���A@0����/#@        ������3@0����/#@        �P^Cy/@��/����?        {�5��(@                z�5��@��/����?        z�5��@                        ��/����?        ��#��@E�JԮD!@        ��#��@                        D�JԮD!@        �P^Cy/@                ���>��,@0����/@0#0# @�k(��"@�cp>@0#0#@��#���?        H�4H�4@��#���?                                H�4H�4@��#�� @�cp>@0#0#�?        �cp>@        ��#�� @        0#0#�?��#�� @                                0#0#�?;��,��@��/����?0#0#@                0#0#@;��,��@��/����?        ;��,��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        z�5��@                        ��/����?        �#���I@���-��*@        6��tSH@���-��@        ���>��,@���-��@        ZLg1��&@                z�5��@���-��@        z�5��@��/����?                ��/����?        z�5��@                        �cp>@        Ey�5A@                z�5��@���-��@        ��#�� @                ��#���?���-��@                ��/���@        ��#���?�cp>@                �cp>@        ��#���?                ���>��@$jW�v%4@��+��+$@��#��@&jW�v%4@��+��+$@��#��@:l��F:2@        ��#�� @9l��F:2@        ��#�� @�cp>@        ��#�� @��/���@                ��/���@        ��#�� @                        ��/����?                ��On�(@        ��#�� @                        ��/����?��+��+$@        ��/����?                ��/����?��+��+$@        ��/����?                        ��+��+$@z�5��@                                H�4H�4@��#��0@��h
�G@,��+��N@<��,��$@鰑5@0#0#�?<��,��$@��/���@        ;��,��@��/���@        ;��,��@��/����?                ��/����?        ;��,��@                        �cp>@        ;��,��@                        E�JԮD1@0#0#�?        ��/���.@                ��/����?0#0#�?        ��/����?                        0#0#�?z�5��@�cp>�9@�A�AN@z�5��@�cp>�9@Y��Y��H@��#�� @D�JԮD1@#0#0F@��#�� @E�JԮD1@�C=�C=<@��#�� @�cp>'@�C=�C=<@��#�� @�cp>'@�C=�C=@��#�� @�cp>'@H�4H�4@��#�� @�cp>@H�4H�4@��#�� @��/����?H�4H�4@        ��/����?H�4H�4@        ��/����?                        H�4H�4@��#�� @��/����?                ��/����?        ��#�� @                        ��/���@                �cp>@                        0#0#@                ��-��-5@                0#0# @                ��)��)3@        �cp>@                ��/����?                ��/���@                        0#0#0@                H�4H�4@                ��8��8*@��#��@D�JԮD!@��+��+@��#��@��/���@��+��+@��#��@��/���@        ��#��@                        ��/���@                        ��+��+@        0����/@                        #0#0&@                0#0# @                vb'vb'"@+�����;@<l��F:B@��+��+T@*�����;@��|��<@H�4H�4(@��b:��*@                ���>��,@��|��<@H�4H�4(@���>��,@鰑%@vb'vb'"@��#�� @/����/#@0#0#@z�5��@E�JԮD!@        ��#�� @E�JԮD!@        ��#�� @                        D�JԮD!@        ��#���?                ;��,��@��/����?0#0#@;��,��@                        ��/����?0#0#@        ��/����?0#0# @                0#0# @        ��/����?                        0#0# @z�5��@��/����?��+��+@z�5��@��/����?0#0#�?z�5��@��/����?        z�5��@                        ��/����?                        0#0#�?                0#0#@        9l��F:2@H�4H�4@        ;l��F:2@0#0#�?        ��/���.@                �cp>@0#0#�?                0#0#�?        �cp>@                ��/����?                ��/����?                        0#0# @        ��/���@V2%S2%Q@        ���-��@�;�;;@        0����/@�;�;;@        ��/���@vb'vb'"@        ��/���@H�4H�4@                H�4H�4@        ��/���@                        H�4H�4@        ��/����?vb'vb'2@        ��/����?0#0# @        ��/����?                        0#0# @                0#0#0@        ��/����?                ��/����?�ڬ�ڬD@                �A�A>@        ��/����?#0#0&@        ��/����?                        #0#0&@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�-#hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKх�h��B�-         �                 ��@s?����T�?$      ��Z�}}@       �                 `m�?�f�Y�c�?�       �a&��xw@       4                 �l�}?�Œ��V�?�       ����VLr@       !                 ��ǻ?��a����?K       y�:�8]@                        @�W?n=:�BY�?.       �J�S@       	                 �"R?�`@s'��?
       �[�_4@                        С=?      �<       ��On�(@������������������������       �               ��/����?������������������������       �               �cp>'@
                        x�8a?>ǵ3���?       �q�ͨ�@������������������������       �               z�5��@������������������������       �               0����/@                        ���@?��~kK��?$       �����K@                         L��?JF�X��?       G�� T�H@                        HR	 ?0#����?       x�߄�C@������������������������       �               �k(��"@                        ��??�N,u��?       ��u�=@������������������������       �      ��	       ������3@                         ���?�Z�	7�?       i~���$@                         ��%?\����?       Q	K��@������������������������       �               ��/����?������������������������       �      �<       z�5��@������������������������       �      ȼ       �cp>@                        ��h�>���/��?       5��o��#@������������������������       �               �cp>@                        ��?�_�A�?       炵�e`@������������������������       �               ��#��@                       �I��F?`%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?                         �$I�?      �<       ���-��@������������������������       �               �cp>@������������������������       �               ��/���@"       +                 �U���xd�$���?       �T�fD@#       *                    �?��?       ��l}�'*@$       %                 �C8�?���Ѯ�?	       ��GQ&@������������������������       �      �<       z�5��@&       '                 �z�?
4=�%�?       �(J��@������������������������       �               ��/����?(       )                 `�z?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      м       ��/����?,       -                 `R|7?h�j���?       \��\�;@������������������������       �      ȼ
       ��b:��*@.       3                  P�"�?�B���?       F��,�,@/       2                 @�K�?Zn����?       ~��Y-"@0       1                  �.�?4=�%�?       �(J��@������������������������       �               ��#�� @������������������������       �               �cp>@������������������������       �               ��#��@������������������������       �               ;��,��@5       �                  8��?�~�fn�?j       zO6�9�e@6       O                  �_�?�#����?h       ^����:e@7       F                 ���`?��J(�?       �nB@8       9                   ��?<
��[,�?       �)�Yj(8@������������������������       �               鰑%@:       ?                 ���?&:�u���?       �j7"�5+@;       >                 ��C�?�`@s'��?       Ei_y,*@<       =                 ��=�?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��/���@@       E                 P
�?��[����?       Hl�_A@A       D                 `s5�?�֪u�_�?       ��?�8@B       C                 0�M�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               �cp>@������������������������       �               0#0#�?G       N                  `s�?���_��?       w@���,(@H       I                 `�?H��aB��?       ����"@������������������������       �               ;��,��@J       K                %I�~�?�@G���?       hu��@������������������������       �               ��/����?L       M                 *\?~�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               H�4H�4@P       {                  �j?H�B����?Q       2&��`@Q       v                 `A��?5�>u��?1       G#l���T@R       o                 P�?�.�j`�?-       ��x�ZS@S       Z                 PRݥ?� ���?       �j?B�qI@T       Y                 ���x?nP�D�?
       �A��P?4@U       V                 ����?H���'0�?	       �C�� T2@������������������������       �               ��/����?W       X                  ��3�?|�6L�n�?       �E#��h0@������������������������       �               ��/����?������������������������       �               ���>��,@������������������������       �      м       ��/����?[       l                 `��?����cY�?       �����>@\       _                   ��?�۫5�?       ��8B!�;@]       ^                  ��g�?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#��@`       c                 �Q+�?�}��	�?       �q�Zz5@a       b                  �}?��F���?       :�.�-'@������������������������       �               鰑%@������������������������       �      �<       ��#���?d       k                  q>�?vutee�?       Q9��#@e       h                 �扨?�� ��?       rp� k@f       g                 �꺖?|��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?i       j                �I�s?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               0#0#@m       n                  pS��?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ��#�� @p       q                 ��L�?���&���?       ���[��:@������������������������       �               ZLg1��&@r       s                  �u��?^n����?       Ӏh��K.@������������������������       �               �cp>@t       u                 PԵ?�����?       �O��(@������������������������       �               <��,��$@������������������������       �      ȼ       ��/����?w       x                 ����?�D�-,�?       �D'ŰO@������������������������       �               0#0#@y       z                ��O�y?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?|       �                 ��.�?"3bc��?        ܁X��
I@}       ~                 �:W>?���=��?       XXs:JB@������������������������       �               ���-��@       �                 H��?躇q@��?       �7t��=@�       �                 �7\?`�s���?       ����'�7@�       �                 (�q?����A�?
       ��]���/@������������������������       �               z�5��@�       �                 �jE?���k�L�?       sk��#@�       �                 x}H�?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 `��?�`@s'��?       Ei_y,*@�       �                 x��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               0����/@������������������������       �      �<       ��/���@�       �                 �ה?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ;��,��@�       �                  Ʒ�?0e��}�?	       ��Se+@������������������������       �      �<       ��On�(@������������������������       �      ܼ       ��#���?������������������������       �      �       H�4H�4@�       �                 @��8?bq�d6�?1       ��u�^�T@�       �                 �%�? ���4w�?        "X��[�L@�       �                 �!�?r]��?       �G��>E@�       �                 ���?���,��?       �>�A@������������������������       �               ��#��@�       �                 p`q�?.����?       ?�:���>@������������������������       �               #0#0&@�       �                 @r��?9�����?
       ��"~��3@������������������������       �               0����/@�       �                 0��?0HA��]�?       ��Ƣ�.@�       �                 ����?Ȕfm���?       ��Z�N@������������������������       �               ��#���?������������������������       �               �cp>@������������������������       �               #0#0&@�       �                 �R�0?<�b���?       �GXvƒ@�       �                 `�N�?�����?       �O��@�       �                 ��>?`n����?       � ��w<@�       �                  s��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               ��#���?������������������������       �      ��       z�5��@������������������������       �               0#0#�?�       �                 �Z��?P��(v��?       �A�s(.@�       �                 �Э�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               ��8��8*@�       �                 ���?�L����?       S2��Â9@������������������������       �               H�4H�4@�       �                  `jS�?�>v�xW�?       行}3|6@�       �                  
N�?\O���?       ��o0@������������������������       �      ��	       鰑%@�       �                 ;��?��íxq�?       %2��-�@�       �                   ���?���mf�?       毠�?b@������������������������       �               0#0#�?������������������������       �      �<       ��/���@������������������������       �               ��#���?������������������������       �               H�4H�4@�       �                 �2��?�d�����?>       \��X@������������������������       �               vb'vb'B@�       �                  �8�?Hy��]0�?)       8.��N@�       �                 0�?�^�F�M�?       ��ޚ�F@�       �                 P��?|�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @�       �                  ��?`,�#6?�?       ���*D@������������������������       �               �;�;;@�       �                 P��?�N�+�?
       ����*@�       �                 �闾?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               ��+��+$@�       �                 Pα�?�~�&��?
       @�]��/@�       �                 �j��?�@G���?       hu��@������������������������       �               0#0#�?�       �                 P���?�;�a
=�?       ��l��@������������������������       �               �cp>@������������������������       �               0#0#�?�       �                  �Ԧ�?      �<       0#0# @������������������������       �               0#0# @������������������������       �               H�4H�4@�t�bh�hhK ��h��R�(KK�KK��h �B�  y�YLGc@�ڕ�]�c@�6k�6�c@y�YLGc@��e�_�b@wb'vb'R@������a@'����-_@k�6k�69@g:��,&S@'jW�v%D@        �k(���E@On��O@@        z�5��@D�JԮD1@                ��On�(@                ��/����?                �cp>'@        z�5��@0����/@        z�5��@                        0����/@        ��k(/D@��/���.@        ��k(/D@D�JԮD!@        ��,���A@��/���@        �k(��"@                �#���9@��/���@        ������3@                z�5��@��/���@        z�5��@��/����?                ��/����?        z�5��@                        �cp>@        ;��,��@0����/@                �cp>@        ;��,��@��/����?        ��#��@                ��#���?��/����?        ��#���?                        ��/����?                ���-��@                �cp>@                ��/���@        ��#��@@��/���@        ��#�� @0����/@        ��#�� @�cp>@        z�5��@                ��#�� @�cp>@                ��/����?        ��#�� @��/����?        ��#�� @                        ��/����?                ��/����?        |�5��8@�cp>@        ��b:��*@                ZLg1��&@�cp>@        z�5��@�cp>@        ��#�� @�cp>@        ��#�� @                        �cp>@        ��#��@                ;��,��@                ��#��P@鰑U@k�6k�69@��#��P@鰑U@��)��)3@z�5��@�e�_��7@H�4H�4@��#���?鰑5@0#0# @        鰑%@        ��#���?鰑%@0#0# @��#���?�cp>@        ��#���?��/����?        ��#���?                        ��/����?                ��/���@                0����/@0#0# @        0����/@0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                �cp>@                        0#0#�?;��,��@�cp>@0#0#@;��,��@�cp>@0#0#�?;��,��@                        �cp>@0#0#�?        ��/����?                ��/����?0#0#�?        ��/����?                        0#0#�?                H�4H�4@Lp�}N@<��18N@��8��8*@]Lg1��F@���-��:@#0#0&@�GpAF@���-��:@H�4H�4@[Lg1��6@h
��6@H�4H�4@���>��,@�cp>@        ���>��,@��/���@                ��/����?        ���>��,@��/����?                ��/����?        ���>��,@                        ��/����?        ��#�� @On��O0@H�4H�4@;��,��@On��O0@H�4H�4@��#��@��/����?                ��/����?        ��#��@                ��#���?��|��,@H�4H�4@��#���?鰑%@                鰑%@        ��#���?                        ��/���@H�4H�4@        ��/���@0#0# @        ��/����?0#0# @                0#0# @        ��/����?                �cp>@                ��/����?                ��/����?                        0#0#@z�5��@                ��#���?                ��#�� @                �k(���5@0����/@        ZLg1��&@                ;��,��$@0����/@                �cp>@        ;��,��$@��/����?        <��,��$@                        ��/����?        ��#���?        ��+��+@                0#0#@��#���?        0#0#�?��#���?                                0#0#�?���>��,@�-����@@0#0# @��b:��*@鰑5@0#0# @        ���-��@        ��b:��*@��|��,@0#0# @���>��@��|��,@0#0# @���>��@���-��@0#0# @z�5��@                ��#���?���-��@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @��#���?�cp>@        ��#���?��/����?                ��/����?        ��#���?                        0����/@                ��/���@        z�5��@                ��#���?                ;��,��@                ��#���?��On�(@                ��On�(@        ��#���?                                H�4H�4@\Lg1��&@�e�_��7@7k�6k�G@<��,��$@/����/#@�z��z�B@<��,��$@D�JԮD!@%S2%S27@;��,��@��/���@#0#06@��#��@                ��#���?��/���@#0#06@                #0#0&@��#���?��/���@#0#0&@        0����/@        ��#���?�cp>@#0#0&@��#���?�cp>@        ��#���?                        �cp>@                        #0#0&@;��,��@��/����?0#0#�?;��,��@��/����?        ��#�� @��/����?        ��#���?��/����?                ��/����?        ��#���?                ��#���?                z�5��@                                0#0#�?        ��/����?�C=�C=,@        ��/����?0#0#�?        ��/����?                        0#0#�?                ��8��8*@��#���?��|��,@��+��+$@                H�4H�4@��#���?��|��,@�C=�C=@��#���?��|��,@0#0#�?        鰑%@        ��#���?��/���@0#0#�?        ��/���@0#0#�?                0#0#�?        ��/���@        ��#���?                                H�4H�4@        /����/#@�
��
�U@                vb'vb'B@        0����/#@n�6k�6I@        ��/���@��+��+D@        ��/����?0#0# @        ��/����?                        0#0# @        ��/����?��)��)C@                �;�;;@        ��/����?#0#0&@        ��/����?0#0#�?                0#0#�?        ��/����?                        ��+��+$@        �cp>@��+��+$@        �cp>@0#0# @                0#0#�?        �cp>@0#0#�?        �cp>@                        0#0#�?                0#0# @                0#0# @                H�4H�4@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ5�;5hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKh��BH4         �                 0�"]?Р��_J�?&      ���}@       �                 0���?7�e���?�       �jXo*4v@       �                 ��C?�&���?�       Tr�G�r@       �                  e�?PZG�g=�?�       ��1��l@       :                 ��*g?�`��Rz�?�       �a&��k@                        ��g^?�/d�-�?<       �ZD�{�Y@                        `%�7? ?�Q���?       ���9@                         �P��?"ذD���?       ������6@	       
                 0��>�f%j��?       ��ꁞ9,@������������������������       �               �cp>@                        @.��>��t� �?       ����x&@������������������������       �               ;��,��@                        �2�Y?\n����?       � ��w<@                        @F��d�$���?       �T�f@                       ��c�@?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ��       z�5��@������������������������       �      ȼ       ��/����?                        `���>lQ��?       �s�=�!@������������������������       �               ��#���?                         _�
?h�r{��?       e�6� @                        �?9?f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �      ��       0����/@                        Ѕ ?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?       '                 ��$?d�އQ�?-       Շ(�fS@       "                 �\͵?��k\��?       nG�
 B@        !                 H,��>      �<
       ��,���1@������������������������       �               ��#��@������������������������       �        	       ��b:��*@#       &                 ��h�>�����?       M��o�g2@$       %                 �P�?���/��?       @z$S��@������������������������       �               �cp>@������������������������       �               z�5��@������������������������       �               z�5��(@(       )                  �Ԧ�?�1�T7;�?       �bF��D@������������������������       �               ��/����?*       7                  ��"?�o����?       ���V��C@+       ,                 �ј<?���M��?       ��� 7@������������������������       �               0����/@-       4                 x�� ?H���'0�?       �C�� T2@.       1                   ��?Hk� ѽ?       �����.@/       0                 h��p?      �<	       ��b:��*@������������������������       �               ��#���?������������������������       �               z�5��(@2       3                 p��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?5       6                    �?      �<       �cp>@������������������������       �               ��/����?������������������������       �               ��/����?8       9                 ~`��      �<
       ��#��0@������������������������       �               ��#�� @������������������������       �               ���>��,@;       h                 �
o?T1e���?P       �+��D]@<       c                 .25Q?xB���t�?(       �e@ǳ�K@=       L                  �Q�?���w�0�?#       kx8nQH@>       K                 (�j5?"�"tb��?       %;���/@?       J                  pjS�?h�H`e��?
       P?��v,@@       A                 �`z?ث���?	       zCOD(@������������������������       �               ��#���?B       I                  ���?�(^:�w�?       Z�� 2&@C       D                 =͗?ھ�R���?       ;�S) $@������������������������       �               0#0#@E       H                 |���?��]ۀ��?       E���O@F       G                 �U�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �               0#0#@������������������������       �      �<       ��#���?������������������������       �      ȼ       ��/����?������������������������       �      м       ��/����?M       T                 pN]�?�����I�?       ��M�8U@@N       S                  ;��?��^���?       ���w!@O       P                    �?xLU���?       h�ҹ^�@������������������������       �               0����/@Q       R                 �r�|?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               0#0#�?U       X                   ��?���/��?       @z$S��7@V       W                 ��Z�?\����?       P	K��@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?Y       b                   +Y�?��߭Q��?       �QVl�0@Z       ]                 PS�?    ���?	       ,x�1�)@[       \                  ���?l@ȱ��?       nm���S@������������������������       �      ��       0����/@������������������������       �               ��#���?^       _                  �g<�?�_�A�?       肵�e`@������������������������       �               ��#��@`       a                 ���?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��/���@d       g                 ���?�`@s'��?       Fi_y,*@e       f                 >�r?      �<       �cp>@������������������������       �               ��/����?������������������������       �               0����/@������������������������       �               ��#���?i       j                 `��?�o���w�?(       ���N@������������������������       �               �cp>@k       n                  ����?:�d��?&       ��ʕbM@l       m                    �?��|��?       ���ĺw@������������������������       �               ��#�� @������������������������       �               0����/@o       t                 `��?$��ʀ�?"       r��I@p       q                 �2*�?�=�Sο?
       ����,@������������������������       �               z�5��(@r       s                 `#p�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?u       v                   E(�?(���� �?       ��ӫo�B@������������������������       �               ��#�� @w       |                  �~��?l8����?       l?�E5=@x       y                 8�K�?�� ��?       rp� k@������������������������       �               ��/���@z       {                 ����?      �<       0#0# @������������������������       �               0#0#�?������������������������       �               0#0#�?}       �                  ���?
Xb���?       N�EBCZ7@~                        P>J�?����X��?	       '��֞&@������������������������       �               ��/����?������������������������       �      �<       ;��,��$@�       �                 x�Gs?��<��?       u=�x�(@������������������������       �               ��/����?�       �                 @��?nP�D�?       �A��P?$@�       �                  �E�?��6L�n�?       �E#��h @������������������������       �               ��/����?������������������������       �      �<       ���>��@������������������������       �      ȼ       ��/����?�       �                 �vQ?f�G���?       �֔�Э#@�       �                 p��!?�~�&��?       ?�]��@�       �                 ���?z�G���?       '5L�`�@������������������������       �               H�4H�4@������������������������       �               �cp>@������������������������       �               0#0# @������������������������       �               ��/����?�       �                 ���\?� ��?!       XP/uM@������������������������       �               z�5��@�       �                 `��?��e�vg�?       ���1��K@�       �                 �yQ?��k~S�?       �2^I�~@@�       �                  ��I? �*�'�?       J���ׅ2@������������������������       �               ��/���@�       �                  ��?��Ñp��?       <7��0�%@������������������������       �               �cp>@�       �                 H8��?����|e�?       �z �B�@�       �                 n�
Q?`�ih�<�?       ��
@�       �                 �-�?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               0#0#@������������������������       �      ȼ       ��/����?�       �                    �?��&���?	       ��G2��,@�       �                ��?d�r{��?       e�6� @�       �                 p��U?�`@s'��?       Ei_y,*@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               ��/����?������������������������       �               ���-��@�       �                 �+�?*ذD���?
       ������6@�       �                 0I��?*��d��?       ��4^$1@�       �                 P`s�?B&Μ�!�?       D3�\r.@������������������������       �               ��/���@������������������������       �               ZLg1��&@������������������������       �      м       ��/����?�       �                    �?      �<       �cp>@������������������������       �               ��/���@������������������������       �               ��/����?�       �                 |�L?�μ���?*       $��~P@�       �                 Ц��?��p�?       ����>?@������������������������       �               �cp>@�       �                    �?����"�?       C��v7<@�       �                  ;��?r^�(���?       � K�h @������������������������       �               0#0#@�       �                 `t��?�3`���?       .�r��@�       �                 ��ɯ?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 ��N�?      �<       0#0# @������������������������       �               0#0#�?������������������������       �               0#0#�?������������������������       �               ��+��+4@�       �                 ��N�?V֡9�2�?       G�8�pA@�       �                 ���?�J�A���?	       3����)@�       �                  p��?�}/W�?       �r�.�%@�       �                 ���!?��^���?       ���w!@������������������������       �               ���-��@������������������������       �               0#0# @������������������������       �               0#0# @������������������������       �               0#0# @�       �                 0�F�?��3�w^�?       /�P�6@�       �                  �Q�?��V���?	       �0��M0@�       �                 p[͔?H[�Jg�?       X�S0f�*@�       �                    �?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?������������������������       �      �<       ;��,��$@������������������������       �               H�4H�4@�       �                  ����?�֪u�_�?       ��?�8@������������������������       �               �cp>@�       �                  ���?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                  �g<�?pό�=�?J       /q�V6b]@�       �                 ���?��h����?       ��[�/@������������������������       �               ��/���@�       �                 P���?v=���?	       � ��R(@������������������������       �               �C=�C=@�       �                 �oW�?�@����?       ���a�@������������������������       �               0#0#@������������������������       �      ȼ       ��/����?�       �                 �L��?�$ ��?>       �34iY@�       �                 `�/c?�a��l�?<       R��B�X@�       �                 �n�?���!��?       �@��&@�       �                 ȃ�?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               ��+��+@�       �                 ��c�?��}n Ӯ?8       G�s��(W@�       �                 p�5i?      �<&       T��N��O@������������������������       �               0#0#�?������������������������       �        %       @�C=�CO@�       �                 �|'�?�ɮ����?       n`E\�=@�       �                 �=�?���};��?       ��;̑�%@������������������������       �               ��+��+@�       �                 �|E�?x�G���?       '5L�`�@������������������������       �               ��/����?�       �                 ����?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@������������������������       �               vb'vb'2@�       �                 �?#�?D�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�t�b�     h�hhK ��h��R�(KK�KK��h �Bh  ��k(/d@z����a@�fm�f�d@�>��d@�-����`@�A�AN@�k(��b@?�)�B]@%S2%S27@�5�װ`@i
���S@S2%S2%1@�5�װ`@�+Q��R@H�4H�4(@B����R@�a#6�;@        ZLg1��&@��|��,@        [Lg1��&@�cp>'@        �k(��"@0����/@                �cp>@        �k(��"@��/����?        ;��,��@                ��#��@��/����?        ��#��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        z�5��@                        ��/����?        ��#�� @���-��@        ��#���?                ��#���?���-��@        ��#���?��/����?                ��/����?        ��#���?                        0����/@                �cp>@                ��/����?                ��/����?        ���b:P@���-��*@        ��#��@@�cp>@        ��,���1@                ��#��@                ��b:��*@                �P^Cy/@�cp>@        z�5��@�cp>@                �cp>@        z�5��@                z�5��(@                �P^Cy?@鰑%@                ��/����?        �P^Cy?@E�JԮD!@        ���>��,@E�JԮD!@                0����/@        ���>��,@��/���@        ���>��,@��/����?        ��b:��*@                ��#���?                z�5��(@                ��#���?��/����?                ��/����?        ��#���?                        �cp>@                ��/����?                ��/����?        ��#��0@                ��#�� @                ���>��,@                ���>��L@��h
�G@H�4H�4(@��#��0@��|��<@��+��+$@�P^Cy/@�cp>7@��+��+$@z�5��@0����/@0#0# @z�5��@�cp>@0#0# @z�5��@��/����?0#0# @��#���?                ��#�� @��/����?0#0# @��#���?��/����?0#0# @                0#0#@��#���?��/����?0#0#@��#���?��/����?                ��/����?        ��#���?                                0#0#@��#���?                        ��/����?                ��/����?        |�5��(@:l��F:2@0#0# @        ���-��@0#0# @        ���-��@0#0#�?        0����/@                ��/����?0#0#�?                0#0#�?        ��/����?                        0#0#�?z�5��(@�cp>'@        z�5��@��/����?        z�5��@                        ��/����?        z�5��@鰑%@        z�5��@���-��@        ��#���?0����/@                0����/@        ��#���?                ;��,��@��/����?        ��#��@                ��#���?��/����?        ��#���?                        ��/����?                ��/���@        ��#���?�cp>@                �cp>@                ��/����?                0����/@        ��#���?                =��,��D@:l��F:2@0#0# @        �cp>@        =��,��D@��/���.@0#0# @��#�� @0����/@        ��#�� @                        0����/@        ������C@鰑%@0#0# @��b:��*@��/����?        z�5��(@                ��#���?��/����?        ��#���?                        ��/����?        �#���9@0����/#@0#0# @��#�� @                ��,���1@0����/#@0#0# @        ��/���@0#0# @        ��/���@                        0#0# @                0#0#�?                0#0#�?��,���1@�cp>@        ;��,��$@��/����?                ��/����?        ;��,��$@                ���>��@0����/@                ��/����?        ���>��@�cp>@        ���>��@��/����?                ��/����?        ���>��@                        ��/����?                0����/@��+��+@        �cp>@��+��+@        �cp>@H�4H�4@                H�4H�4@        �cp>@                        0#0# @        ��/����?        �P^Cy/@�+Q��B@H�4H�4@z�5��@                z�5��(@�+Q��B@H�4H�4@��#���?�cp>�9@H�4H�4@        ��On�(@H�4H�4@        ��/���@                0����/@H�4H�4@        �cp>@                ��/����?H�4H�4@        ��/����?H�4H�4@        ��/����?0#0# @        ��/����?                        0#0# @                0#0#@        ��/����?        ��#���?���-��*@        ��#���?���-��@        ��#���?�cp>@                �cp>@        ��#���?                        ��/����?                ���-��@        ZLg1��&@�cp>'@        [Lg1��&@�cp>@        ZLg1��&@��/���@                ��/���@        ZLg1��&@                        ��/����?                �cp>@                ��/���@                ��/����?        [Lg1��&@E�JԮD1@�z��z�B@��#���?��/���@��8��8:@        �cp>@        ��#���?��/����?��8��8:@��#���?��/����?H�4H�4@                0#0#@��#���?��/����?0#0# @��#���?��/����?                ��/����?        ��#���?                                0#0# @                0#0#�?                0#0#�?                ��+��+4@<��,��$@���-��*@#0#0&@        ���-��@H�4H�4@        ���-��@0#0#@        ���-��@0#0# @        ���-��@                        0#0# @                0#0# @                0#0# @;��,��$@���-��@��+��+@<��,��$@��/����?0#0#@;��,��$@��/����?0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?;��,��$@                                H�4H�4@        0����/@0#0#�?        �cp>@                ��/����?0#0#�?                0#0#�?        ��/����?        ��#���?0����/#@������Z@        0����/@#0#0&@        ��/���@                ��/����?#0#0&@                �C=�C=@        ��/����?0#0#@                0#0#@        ��/����?        ��#���?0����/@D�s?��W@��#���?��/���@<k�6k�W@��#���?��/����?��+��+@��#���?��/����?        ��#���?                        ��/����?                        ��+��+@        �cp>@��
�pV@                T��N��O@                0#0#�?                @�C=�CO@        �cp>@��8��8:@        �cp>@0#0# @                ��+��+@        �cp>@H�4H�4@        ��/����?                ��/����?H�4H�4@        ��/����?                        H�4H�4@                vb'vb'2@        ��/����?0#0#�?        ��/����?                        0#0#�?�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJi4�hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KKم�h��Bx/         �                  t0�?07�LJ�?      �8��Gs}@       y                 ����?�% ooV�?�       v+8���u@       @                 @ۣ?��l�.�?�       ��ߏ�p@       +                 ���@?����?_       �mtL�	d@                        @�W?f��4�?H       1�s��\@                         �{��?�3�g�?       ׵5��2@       
                  q�?�(�����?       ��0��0@       	                 @���>���/��?       @z$S��@������������������������       �               �cp>@������������������������       �               z�5��@                        @Ws�?�^�#΀�?	       N�{��A%@������������������������       �      ��       D�JԮD!@                        hì+?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ܼ       ��#�� @                        �����6�	lw�?;       �2�xQX@                        �_?�����?       ��/̸IC@                        �ìW?����5�?       B�)�B=@������������������������       �               ��/���@                        ���g?�:�^���?       ��]�ڕ5@������������������������       �               z�5��(@                        p�j?L���'0�?       �C�� T"@������������������������       �               ��/����?                        0vb�?��6L�n�?       �E#��h @                        �j��?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               z�5��@������������������������       �               �k(��"@       (                  �u��?�g	9�H�?!       �<5�8YM@        '                ���1�?���/��?       @z$S��@!       $                  �q�?����?       ��X�)B@"       #                 �a{?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?%       &                 L�5E?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?������������������������       �      �<       ��/����?)       *                 P>_�? С�K�?       ��Я[[J@������������������������       �               �#���I@������������������������       �      �<       ��/����?,       -                  `��?P-zl��?       2]�p�-F@������������������������       �               ��#��@.       9                 ����?f9��;3�?       �ll�D@/       8                    �?P?�腷�?       4֖v�<@0       5                  �Q�?F��3��?       �_q>c3@1       4                 ��c?�0�~��?	       r��GQ1@2       3                �-~�?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �               ���-��*@6       7                 �Z�?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?������������������������       �               E�JԮD!@:       ?                    �?�����?       �Ä�>c(@;       >                  ����?��t� �?       ����x&@<       =                 Ĉ�{?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ��       ���>��@������������������������       �      м       ��/����?A       j                  ���?~��<w6�?:       ����V*[@B       ]                 0vb�?�u�!��?)       �	RؘYR@C       L                 �5W�?k�<	N��?       ����E@D       G                  �P�?:��?�D�?       �\��(�%@E       F                   .p�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?H       I                 hU�<?h����?       �����!@������������������������       �               0#0#@J       K                 ����?hutee�?       Q9��@������������������������       �               ��/����?������������������������       �               H�4H�4@M       R                 \F�M?ҭ�8&S�?       �x��T&?@N       Q                  @?��?@��~d��?       7E���*@O       P                 @�C�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �      ��       鰑%@S       \                  Ւ?�C>�?       �1�m�1@T       [                 ��f?(��5�?       ��~���%@U       V                 P,��?2�c3���?       �uk��!@������������������������       �               ��#�� @W       X                  �P�?��|��?       ���ĺw@������������������������       �               ��/���@Y       Z                 �΅�?^n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               0#0# @������������������������       �               ���-��@^       g                  �E�?�p5Z4�?       � .J�F?@_       d                 `���?�5��E��?       �Ȍ�p;@`       c                 Pk�?���q���?       �:-ߩ�+@a       b                  �\�?�@G���?       hu��@������������������������       �               0#0# @������������������������       �               �cp>@������������������������       �               z�5��@e       f                 0�� ?      �<       ��b:��*@������������������������       �               ;��,��@������������������������       �               ��#�� @h       i                    �?      �<       ��/���@������������������������       �               �cp>@������������������������       �               ��/����?k       r                 ��L�?`��ʸ��?       P�
|�A@l       m                 �9��?���q���?       �:-ߩ�@������������������������       �               ��#�� @n       o                 n�
Q?����]L�?       N66�ͯ@������������������������       �               �cp>@p       q                 L��?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?s       v                  +�?l<
H<�?       �J�E<@t       u                 MԦ?�|2N��?       �3K}@������������������������       �               z�5��@������������������������       �               0#0# @w       x                  @���?@4�+W�?
       ����%7@������������������������       �      ��	       #0#06@������������������������       �      �<       ��/����?z       �                 �6Sz?�F��1��?7       �K �*�T@{       �                 �\��?�8�E��?(       O+A2FP@|       �                  8��?�^�D�?!       TIo-��J@}       �                 P���?��Rb���?       3m
��I@~       �                  �x��?�m�=�k�?       j���G@       �                 ��jm?      �<       �e�_��7@������������������������       �               ��On�(@������������������������       �               �cp>'@�       �                   �P�?�<=��c�?       0ne��Y7@������������������������       �               ��#�� @�       �                 ��Ĳ?�}>D�P�?       �狢G5@�       �                 Pd�?�Ș���?       �̨	�>4@������������������������       �               0#0#�?�       �                   �0�?�����o�?       ]���v<3@�       �                 Z��?���mf�?       毠�?b@������������������������       �               0#0#�?������������������������       �      �<       ��/���@������������������������       �               ��|��,@������������������������       �      �<       ��#���?�       �                 xQ}�?|�G���?       ��%�|@������������������������       �               0#0# @������������������������       �      �<       ��/����?�       �                 �3ܦ?     ��<       0#0# @������������������������       �               0#0#�?������������������������       �               0#0#�?�       �                 0]��?z�G���?       '5L�`�'@�       �                  PV��?|��`p��?       f;3@��!@������������������������       �               �cp>@������������������������       �      �<       H�4H�4@������������������������       �      Լ       �cp>@�       �                 X���?8��b�?       %�|�1@�       �                 (�œ?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      ��       �A�A.@�       �                 �8��?�-Y�M�?M       �5��^@�       �                 l��t?�!�����?       ��9�H@�       �                 @��8?��J67�?       �J���?@�       �                  ��?�;<`�?       �q�:>7@������������������������       �               ���>��@�       �                    �?_f"��?
        ��Um�/@�       �                 �|��?|(� C�?	       sۋɬ�+@������������������������       �               H�4H�4@�       �                 ��{�?&��5�?       ��~���%@�       �                 0���?���`�?       ��
�Me@�       �                  u��?��n��?       �-H�\@�       �                �E9�?�֪u�_�?       ��?�8@�       �                 4zM�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �               z�5��@������������������������       �               0#0# @�       �                 0��?��^���?       ���w!@������������������������       �               0#0# @������������������������       �               ���-��@�       �                 0��?xr����?
       Qz�i0@������������������������       �               0#0# @�       �                 ���?�v�;B��?       ՟���	 @�       �                 ��?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?������������������������       �               H�4H�4@�       �                 P��m?B+�Y�P�?0       �N�p��Q@�       �                    �?YX�\�?       �˱d�C@�       �                  ��?��[����?       Gl�_A@������������������������       �      ��       0����/@������������������������       �               0#0# @�       �                 pNh�?�����6�?       b�i�8r@@�       �                 � �8?
�x��>�?       �	�{ �9@�       �                 �P�?�78���?       [�i:e2@�       �                  v�?�@G���?       hu��@������������������������       �               ��/����?�       �                 P��?~�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                pn�ǣ?��p\�?       �����J,@������������������������       �        
       H�4H�4(@�       �                 �O׶?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?�       �                 (�A�?3y�d��?       �)h�2@������������������������       �               ��#���?�       �                   ���?�;�a
=�?       ��l��@�       �                 t�N�?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?�       �                 0�c�?      �<       ��/���@������������������������       �               ��/����?������������������������       �               ��/����?������������������������       �               �C=�C=@�       �                 �m۶?      �<       0#0#@@������������������������       �               0#0#@������������������������       �               �C=�C=<@�t�bh�hhK ��h��R�(KK�KK��h �BX  g:��,&c@�H��tXe@~��~�gb@}�5�wa@Y<�œb@D�A�P@Gy�5a@��h
�W@��)��)C@V^CyeZ@���-��J@0#0#�?:��P^�V@�cp>�9@        z�5��@��On�(@        ��#��@��On�(@        z�5��@�cp>@                �cp>@        z�5��@                ��#���?/����/#@                D�JԮD!@        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                bCy��T@���-��*@        ���>��<@0����/#@        ������3@0����/#@                ��/���@        ������3@��/����?        z�5��(@                ���>��@��/����?                ��/����?        ���>��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        z�5��@                �k(��"@                �>��nK@��/���@        z�5��@�cp>@        z�5��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#�� @                ��#���?                ��#���?                        ��/����?        �#���I@��/����?        �#���I@                        ��/����?        �P^Cy/@�a#6�;@0#0#�?��#��@                \Lg1��&@�a#6�;@0#0#�?��#�� @��On�8@0#0#�?��#�� @On��O0@0#0#�?        On��O0@0#0#�?        �cp>@0#0#�?        �cp>@                        0#0#�?        ���-��*@        ��#�� @                ��#���?                ��#���?                        E�JԮD!@        �k(��"@�cp>@        �k(��"@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ���>��@                        ��/����?        �P^Cy?@%jW�v%D@�z��z�B@{�5��8@:l��F:B@H�4H�4(@;��,��@���-��:@��+��+$@��#���?�cp>@�C=�C=@��#���?��/����?                ��/����?        ��#���?                        ��/����?�C=�C=@                0#0#@        ��/����?H�4H�4@        ��/����?                        H�4H�4@��#��@�e�_��7@H�4H�4@        ��On�(@0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                鰑%@        ��#��@�cp>'@0#0# @��#��@0����/@0#0# @��#��@0����/@        ��#�� @                ��#�� @0����/@                ��/���@        ��#�� @��/����?        ��#�� @                        ��/����?                        0#0# @        ���-��@        ������3@0����/#@0#0# @������3@�cp>@0#0# @z�5��@�cp>@0#0# @        �cp>@0#0# @                0#0# @        �cp>@        z�5��@                ��b:��*@                ;��,��@                ��#�� @                        ��/���@                �cp>@                ��/����?        z�5��@��/���@k�6k�69@z�5��@�cp>@0#0#�?��#�� @                ��#���?�cp>@0#0#�?        �cp>@        ��#���?        0#0#�?                0#0#�?��#���?                z�5��@��/����?H�4H�48@z�5��@        0#0# @z�5��@                                0#0# @        ��/����?#0#06@                #0#06@        ��/����?        z�5��@o��F:lI@�C=�C=<@z�5��@��On�H@H�4H�4(@z�5��@h
��F@H�4H�4@z�5��@h
��F@0#0#@z�5��@鰑E@0#0# @        �e�_��7@                ��On�(@                �cp>'@        z�5��@;l��F:2@0#0# @��#�� @                ��#���?:l��F:2@0#0# @        :l��F:2@0#0# @                0#0#�?        :l��F:2@0#0#�?        ��/���@0#0#�?                0#0#�?        ��/���@                ��|��,@        ��#���?                        ��/����?0#0# @                0#0# @        ��/����?                        0#0# @                0#0#�?                0#0#�?        �cp>@H�4H�4@        �cp>@H�4H�4@        �cp>@                        H�4H�4@        �cp>@                ��/����?0#0#0@        ��/����?0#0#�?        ��/����?                        0#0#�?                �A�A.@��b:��*@�cp>�9@��+��+T@[Lg1��&@��On�(@H�4H�48@[Lg1��&@�cp>'@vb'vb'"@ZLg1��&@0����/@�C=�C=@���>��@                ��#��@0����/@�C=�C=@��#��@0����/@��+��+@                H�4H�4@��#��@0����/@0#0# @��#���?0����/@0#0# @��#���?0����/@0#0#�?        0����/@0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?                �cp>@        ��#���?                                0#0#�?z�5��@                                0#0# @        ���-��@0#0# @                0#0# @        ���-��@                ��/����?�A�A.@                0#0# @        ��/����?�C=�C=@        ��/����?0#0#�?                0#0#�?        ��/����?                        H�4H�4@��#�� @���-��*@�C=�C=L@��#�� @���-��*@H�4H�48@        0����/@0#0# @        0����/@                        0#0# @��#�� @D�JԮD!@#0#06@��#�� @D�JԮD!@�A�A.@��#���?�cp>@�C=�C=,@        �cp>@0#0#�?        ��/����?                ��/����?0#0#�?                0#0#�?        ��/����?        ��#���?        ��8��8*@                H�4H�4(@��#���?        0#0#�?��#���?                                0#0#�?��#���?�cp>@0#0#�?��#���?                        �cp>@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/���@                ��/����?                ��/����?                        �C=�C=@                0#0#@@                0#0#@                �C=�C=<@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�ThFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK兔h��B2         �                 �6Sz?����T�?,      ��Z�}}@       g                 0-3�?j�L�S�?�       (,����w@                           �G�?.�n�^�?y       ���Ug@                        �%��?�w��?       
�H�
�G@       
                  ��~�?X-zl��?       3]�p�-F@                        �$�N?F���'0�?       �C�� T"@������������������������       �               z�5��@       	                 @F�f%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?                        �q�3?y>�S��?       F̴9��A@                        Pc��?P�,��?       �t5ë6@                        ,*���\���A�?       .gX\-@                       ��z�? e��}�?
       ��Se+@������������������������       �               ��#���?������������������������       �        	       ��On�(@������������������������       �      �<       ��#���?                         �x?����?       ��X�)B @                        x���?\n����?       � ��w<@                        ��?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?������������������������       �               ��#�� @                        82�?�+�z���?	       LGh��
)@������������������������       �               鰑%@                           �?z�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?                       8�|�?      �<       z�5��@������������������������       �               ��#�� @������������������������       �               ��#���?!       V                 ���@?ܕ���?Z       7�6ga@"       '                 ��V?L����&�?E       �7�Fg�[@#       &                 ��J�?��|��?
       ���ĺw+@$       %                 p�3G?6�c3���?       �uk��!@������������������������       �               ��#��@������������������������       �               0����/@������������������������       �      ȼ       0����/@(       U                  U\�?�����?;       ���o:X@)       <                 P��?���_��?9       ��7³�V@*       5                 ����?P�؈�w�?       q���S#G@+       2                 �Q�?`����?       �Fx�v�5@,       /                 ��p?�hK)�?
       �h��K�2@-       .                  Pmj�?\����?       P	K��@������������������������       �               ��/����?������������������������       �               z�5��@0       1                 ��aӾ      �<       ZLg1��&@������������������������       �               ��#��@������������������������       �               ���>��@3       4                 x#]?b%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?6       ;                  ��d�? ��K��?       ���0�8@7       :                ����.?��6L�n�?       �E#��h @8       9                 .6U@?`n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      �<       ;��,��@������������������������       �      м
       ��#��0@=       >                 �;�b?�YX�io�?       ;³��F@������������������������       �               ��/����??       L                 Ш��?���Ѯ�?       ��GQF@@       G                 �m��?<9�)\e�?       ��)8@A       D                 � 1?�q���?       ��|�^1@B       C                   �x�?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?E       F                  �ޖ?�=�Sο?	       ����,@������������������������       �               ��b:��*@������������������������       �      ȼ       ��/����?H       K                  �JV�?�`@s'��?       Di_y,*@I       J                ���[�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?������������������������       �      ȼ       0����/@M       R                 `���?�3��F��?       nf9t{y4@N       Q                 �.م?Hk� ѽ?
       �����.@O       P                    �?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@������������������������       �      ��       <��,��$@S       T                 ��=�?ܗZ�	7�?       j~���@������������������������       �               ��/����?������������������������       �               z�5��@������������������������       �      �       ��+��+@W       Z                  ����?��Ұ��?       �1��<@X       Y                 Pc	�? ��c`�?
       $��t5)@������������������������       �      ��	       �cp>'@������������������������       �      �<       ��#���?[       \                 XJO
?�A&w(�?       �]��0@������������������������       �               ��/���@]       f                  0p��?����?       �Ä�>c(@^       e                  ���?Xn����?       ��Y-"@_       d                 �w2�?�����?       ��X�)B @`       a                 ����?\����?       P	K��@������������������������       �               ��#��@b       c                  `�J�?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?������������������������       �      м       ��/����?������������������������       �      ȼ       z�5��@h       �                 ��n�?��R�L��?z       �jb��g@i       �                 �x�y?Cr3����?9       ��D
�BV@j       y                    �?b�����?       L��P�B@k       v                 p��!?�dI�Ɲ�?       ɑ�P>z2@l       m                 `��?A��NV=�?       �t�ܲ@������������������������       �               0#0#�?n       o                 �?su? �Z�ܙ�?       c����@������������������������       �               ��#���?p       u                 GW�d?��íxq�?       %2��-�@q       r                 йu�?����]L�?       N66�ͯ@������������������������       �               �cp>@s       t                  Џ~�?�J���?       ��*]Y @������������������������       �               ��#���?������������������������       �               0#0#�?������������������������       �      м       ��/����?w       x                 ���?      �<       鰑%@������������������������       �               ��/����?������������������������       �               D�JԮD!@z       �                   �g�?R����?       �|�c�2@{       |                 ��q?a{���?       �~8�31@������������������������       �               0#0#@}       ~                 �ݯ�?�W�-q�?	       �|_,��)@������������������������       �               �cp>@       �                  P�"�?�g�(�>�?       �F�V;$@�       �                 h�R?���WW�?       �j�S@�       �                 04�?�|2N��?       �3K}@������������������������       �               z�5��@������������������������       �               0#0# @������������������������       �      ȼ       ��/����?������������������������       �               0#0#@������������������������       �      м       ��/����?�       �                 �p�?��X	]�?!       ���+��I@�       �                 T��p?f�B��#�?       J[���5@������������������������       �               �cp>@�       �                 ��?;���Jt�?       j���3@�       �                 �$�?����?
       }�5�1@�       �                 0�{?T����1�?       ��;9�@������������������������       �               0#0# @������������������������       �               ��#��@�       �                 �W��?���};��?       ��;̑�%@������������������������       �               ��/����?�       �                 p�v�?�@����?       ���a�#@������������������������       �               �C=�C=@�       �                 p-3�?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?�       �                 Db?      �<       ��/����?������������������������       �               ��/����?������������������������       �               ��/����?�       �                 p-�?�N,u��?       ��u�=@�       �                 ���}?`n����?       ��Y-"@������������������������       �               ��/����?�       �                 ��{�?d����?       P	K��@������������������������       �               z�5��@������������������������       �      ȼ       ��/����?�       �                 ����?��#�Ѵ�?       �)�B�4@������������������������       �        
       ���>��,@�       �                 ��'�?�����?       �O��@������������������������       �               ��/����?������������������������       �               ;��,��@�       �                  ���?�'���h�?A       _ �$�Y@�       �                 �I�?>�9�6%�?/       �L˜G�R@�       �                  `S��?�|-7�X�?+       d�E�$�Q@�       �                 Џ�B?�^P-C�?&       K����O@�       �                 �ڡ�?T�����?       D�JS,B@�       �                    �?j�ld���?       ���$]Z:@�       �                 ���?��[����?       Hl�_A@������������������������       �               0����/@������������������������       �               0#0# @�       �                  �g<�?$�Zh�=�?	       �"<2�3@�       �                 p���?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@�       �                 ��2�?�QG�u�?       ALx��.@�       �                 0?��,���?       "C�s��,@������������������������       �               ���-��*@������������������������       �               0#0#�?������������������������       �      ܼ       ��#���?�       �                     �?;ʁ���?       ^]*_�#@������������������������       �               ��/����?�       �                 ���?����?       �a�E�$ @�       �                 p�?�D�-,�?       �D'ŰO@�       �                 �C8�?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               0#0#@�       �                 0��?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 �N��?����x�?       �ra6�:@������������������������       �               ��On�8@�       �                 ؗ�j?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?�       �                 h�B?     ��<       �C=�C=@������������������������       �               0#0#@������������������������       �               H�4H�4@�       �                 ��cb?؃���?       ��X�)B@������������������������       �      �<       z�5��@������������������������       �      �<       ��/����?�       �                 pdJ�?�'1n 6�?       E��N:@������������������������       �      ȼ
       �C=�C=,@�       �                 �ڡS?��n?�?       �ZhiX�'@�       �                 �}��?����]L�?       N66�ͯ@�       �                 0Ϯ�?��q�R�?       C}Ԥ@������������������������       �               ��#���?�       �                 �؉�?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                 �lw?X�ih�<�?       ��
@������������������������       �               H�4H�4@������������������������       �      ȼ       ��/����?�       �                 ��;�? G��?9       ���%��W@������������������������       �        #       -��+��N@�       �                 ܆�?�6��b�?       &�|�A@�       �                 �� �?����|e�?       �z �B�@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                  ��^�? �v}�?       ���5>@�       �                 ����?X�ih�<�?       ��
@������������������������       �               ��/����?������������������������       �               H�4H�4@�       �                 ��Q�?      �<       %S2%S27@������������������������       �               0#0# @������������������������       �               ��-��-5@�t�bh�hhK ��h��R�(KK�KK��h �Bx  y�YLGc@�ڕ�]�c@�6k�6�c@y�YLGc@�z����c@8��8�cP@��+[@����Q@H�4H�4@�k(��2@�a#6�;@0#0#�?�P^Cy/@�a#6�;@0#0#�?���>��@��/����?        z�5��@                ��#���?��/����?                ��/����?        ��#���?                ��#�� @�cp>�9@0#0#�?��#�� @��|��,@        ��#�� @��On�(@        ��#���?��On�(@        ��#���?                        ��On�(@        ��#���?                z�5��@��/����?        ��#��@��/����?        ��#��@��/����?        ��#��@                        ��/����?                ��/����?        ��#�� @                        �cp>'@0#0#�?        鰑%@                ��/����?0#0#�?                0#0#�?        ��/����?        z�5��@                ��#�� @                ��#���?                :��P^�V@h
��F@��+��+@�b:���S@�cp>�9@��+��+@��#��@/����/#@        ��#��@0����/@        ��#��@                        0����/@                0����/@        C����R@On��O0@��+��+@B����R@On��O0@        ���#8E@��/���@        �k(��2@�cp>@        ��,���1@��/����?        z�5��@��/����?                ��/����?        z�5��@                ZLg1��&@                ��#��@                ���>��@                ��#���?��/����?                ��/����?        ��#���?                �,����7@��/����?        ���>��@��/����?        ��#�� @��/����?                ��/����?        ��#�� @                ;��,��@                ��#��0@                ��#��@@��On�(@                ��/����?        ��#��@@�cp>'@        �P^Cy/@D�JԮD!@        ���>��,@�cp>@        ��#���?��/����?        ��#���?                        ��/����?        ��b:��*@��/����?        ��b:��*@                        ��/����?        ��#���?�cp>@        ��#���?��/����?                ��/����?        ��#���?                        0����/@        ��,���1@�cp>@        ���>��,@��/����?        ��#��@��/����?                ��/����?        ��#��@                <��,��$@                z�5��@��/����?                ��/����?        z�5��@                                ��+��+@;��,��$@;l��F:2@        ��#���?�cp>'@                �cp>'@        ��#���?                �k(��"@���-��@                ��/���@        �k(��"@�cp>@        z�5��@�cp>@        z�5��@��/����?        z�5��@��/����?        ��#��@                ��#�� @��/����?                ��/����?        ��#�� @                        ��/����?                ��/����?        z�5��@                ]Lg1��F@鰑U@����M@��,���A@�]�ڕ�?@#0#06@;��,��@$jW�v%4@H�4H�4(@��#�� @��|��,@0#0# @��#�� @��/���@0#0# @                0#0#�?��#�� @��/���@0#0#�?��#���?                ��#���?��/���@0#0#�?��#���?�cp>@0#0#�?        �cp>@        ��#���?        0#0#�?��#���?                                0#0#�?        ��/����?                鰑%@                ��/����?                D�JԮD!@        z�5��@�cp>@��+��+$@z�5��@��/���@��+��+$@                0#0#@z�5��@��/���@H�4H�4@        �cp>@        z�5��@��/����?H�4H�4@z�5��@��/����?0#0# @z�5��@        0#0# @z�5��@                                0#0# @        ��/����?                        0#0#@        ��/����?        Lp�}>@�cp>'@��+��+$@��#��@��/���@��+��+$@        �cp>@        ��#��@0����/@��+��+$@��#��@�cp>@��+��+$@��#��@        0#0# @                0#0# @��#��@                        �cp>@0#0# @        ��/����?                ��/����?0#0# @                �C=�C=@        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?                ��/����?                ��/����?        �#���9@��/���@        z�5��@�cp>@                ��/����?        z�5��@��/����?        z�5��@                        ��/����?        ������3@��/����?        ���>��,@                ;��,��@��/����?                ��/����?        ;��,��@                <��,��$@f#6�aJ@�z��z�B@�k(��"@z%jW�vH@0#0#0@z�5��@�e�_��G@0#0#0@z�5��@�e�_��G@vb'vb'"@z�5��@h
��6@0#0# @��#��@0����/3@H�4H�4@        0����/@0#0# @        0����/@                        0#0# @��#��@��|��,@0#0#�?z�5��@��/����?                ��/����?        z�5��@                ��#���?���-��*@0#0#�?        ���-��*@0#0#�?        ���-��*@                        0#0#�?��#���?                ��#�� @�cp>@��+��+@        ��/����?        ��#�� @��/����?��+��+@��#���?        ��+��+@��#���?        0#0#�?                0#0#�?��#���?                                0#0#@��#���?��/����?                ��/����?        ��#���?                        �cp>�9@0#0#�?        ��On�8@                ��/����?0#0#�?        ��/����?                        0#0#�?                �C=�C=@                0#0#@                H�4H�4@z�5��@��/����?        z�5��@                        ��/����?        ��#���?��/���@��-��-5@                �C=�C=,@��#���?��/���@�C=�C=@��#���?�cp>@0#0#�?��#���?��/����?0#0#�?��#���?                        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?                ��/����?H�4H�4@                H�4H�4@        ��/����?                ��/����?2��-�rW@                -��+��N@        ��/����?0#0#@@        ��/����?H�4H�4@        ��/����?                        H�4H�4@        ��/����?�s?�s?=@        ��/����?H�4H�4@        ��/����?                        H�4H�4@                %S2%S27@                0#0# @                ��-��-5@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ5�R/hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK݅�h��BX0         �                  t0�?��%��G�?*      ��m9N�}@       �                 pY7e?�}���3�?�       ��
G�u@       �                  ��?h��t���?�       �ۃ���r@       7                 ��_i? ��acm�?�        ����r@                        �$?Z?��Ս7�?I       ���^�^@                        �y������'��?       �v�9��4@                        ��l?|���A�?
       /gX\-@                        .25Q?e��}�?	       ��Se+@	                        ��IL?�^�#΀�?       O�{��A%@
                        ��B?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �      ��       D�JԮD!@������������������������       �               �cp>@������������������������       �      ܼ       ��#���?                         ����?      �<       z�5��@������������������������       �               ��#�� @������������������������       �               ��#��@       *                 �b)U?�{F���?;       ")g89tY@                        ��$?5��O�?(       <>�\��Q@                        @��>�	�� ��?       ?�x��>@                        @��>�d�$���?       �T�f@������������������������       �               ��#�� @                        �7r?\n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               �#���9@       )                 ��K�?�d�$���?       �T�fD@                        `ۭ1?��Ӭ%�?       ޅ��pC@������������������������       �               �cp>@       (                 `�ռ?��k\��?       nG�
 B@        '                 ��E?l\Cl[��?       >�s�d�9@!       &                 �G�?�B���?       F��,�,@"       %                  �g<�?bn����?       ~��Y-"@#       $                    �?Ĕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?������������������������       �               ;��,��@������������������������       �      ��       ;��,��@������������������������       �      ȼ       \Lg1��&@������������������������       �               <��,��$@������������������������       �      �<       ��/����?+       2                 05�|?kA�7A��?       ��{n�
>@,       1                  �/�?�d�$���?
       <��#�.@-       0                   .p�?X�s�	�?	       f���*@.       /                 �}��?����?       ��X�)B@������������������������       �               ��/����?������������������������       �      ��       z�5��@������������������������       �      м       �k(��"@������������������������       �      ȼ       ��/����?3       6                 `K�?ʂ�O���?	       �O�
|-@4       5                 �ڭ?�}	;	�?       uK�>4%@������������������������       �               0#0#�?������������������������       �      ��       0����/#@������������������������       �               ��#��@8                        P>J�?��"U��?j       ��[t�d@9       \                 ���?��YMP��?F       >��$C)[@:       O                 `��?�0�w�?-       }';�Q@;       <                     �?<a_)��?#       d����J@������������������������       �               ���-��*@=       >                  �\�?*�W��~�?       ����C@������������������������       �               ��#���??       F                  ��?�	/����?       c�NzC@@       E                 �I?�4��v�?       �Y-"�'@A       D                 ��?������?       �4^$4�#@B       C                 ��K?      �<       ���-��@������������������������       �               ��/����?������������������������       �               0����/@������������������������       �      ȼ       z�5��@������������������������       �               ��#�� @G       L                 ��_?���C��?       >W=��;@H       K                 (�Q�? �v���?       )f�n8@I       J                 �G��?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �               h
��6@M       N                 J}P?ln����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @P       Y                 �	I�?Hh��ې�?
       ��Ւ1@Q       R                 �X�}?�_�A�?       肵�e`,@������������������������       �               ;��,��@S       T                 p���?� �_rK�?       J�@��"@������������������������       �               z�5��@U       V                 @�]�?d%@�"�?       ��[�@������������������������       �               ��/���@W       X                 0�2�?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?Z       [                 @�#�?�� ��?       rp� k@������������������������       �               0#0#�?������������������������       �      �<       ��/����?]       p                    �?p���?       X�FCC@^       _                 ��t?0�Cx@��?       X�k�30@������������������������       �               ��/����?`       o                 ��_?�fB��?       �^q�,,@a       l                 0�ߢ?����W�?
       �`���@*@b       k                ��X�p?����?       ���"�X$@c       h                  h�B?�W�w��?       �'DQm"@d       e                 `�г?��ڰ�x�?       �K�f�@������������������������       �               z�5��@f       g                 `0��?T����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @i       j                  .p�?\n����?       � ��w<@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �      ȼ       ��/����?m       n                 ����?Z%@�"�?       ��[�@������������������������       �               ��/����?������������������������       �      �<       ��#���?������������������������       �      м       ��/����?q       ~                 p~�u?�����?       W!��6@r       s                 �p�?ҟ��X�?       l�n�/4@������������������������       �               �C=�C=@t       {                 �s%�?����W�?	       �`���@*@u       z                 .�X?X�j���?       ���z"@v       y                 �-�?��6L�n�?       �E#��h @w       x                 Ш��?`n����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �      �<       ;��,��@������������������������       �      �<       ��#���?|       }                  ���?�@G���?       hu��@������������������������       �               �cp>@������������������������       �               0#0#�?������������������������       �      м       ��/����?�       �                 ���?��5���?$       ̪&K[M@�       �                 �闾?(��j�?       �4Z��H@�       �                 h��1?�3`���?       -�r�� @�       �                 I��?���/��?       V��7�@������������������������       �               ��/����?������������������������       �               ��#�� @������������������������       �               0#0#@�       �                   �0�? ?6��,�?       us���D@�       �                 Pq��?��x�,�?        �z��?@�       �                 ��k?X7uV��?       �l}�'�:@�       �                 ��??���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?�       �                 �-�?      �<       z�5��8@������������������������       �               ��#���?������������������������       �               �,����7@�       �                  �9��?4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @�       �                 �^�?ޗZ�	7�?       j~���$@������������������������       �               ;��,��@�       �                 @���?& k�Lj�?       �q��l}@������������������������       �               ��/����?�       �                    �?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 ���U?[�H�q�?       ��	0�!@�       �                 �(��?�֪u�_�?       ��?�8@������������������������       �               0#0#�?������������������������       �      ��       0����/@�       �                  �6�?�D#���?       �B�j@������������������������       �               ��#���?������������������������       �               0#0# @�       �                 ��I�?�:[��G�?       �O�;�]!@�       �                 �̚y?|�G���?       ��%�|�?������������������������       �               ��/����?������������������������       �               0#0#�?������������������������       �      �<       ���-��@�       �                 ��9�?��ޖ��?$       �3�J@�       �                 @F���-�\�?#       �(gJ@�       �                 �?�?|�G���?       ��%�|@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 0�/�?r����?       �y���!H@�       �                 �\ͥ?      �<       k�6k�69@������������������������       �               0#0#�?������������������������       �               H�4H�48@�       �                 �w��?���q��?       �?8��7@������������������������       �               ��/����?�       �                 ܆�?�^�F�M�?       ��ޚ�6@�       �                 �k�?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                  N��?8L�0�h�?       l�e�3@������������������������       �        
       vb'vb'2@������������������������       �      �<       ��/����?������������������������       �      �<       ��/����?�       �                   ҏ�?Z�4-���?M       �G�8^@�       �                 0I��?�֪u�_�?       ��?�8'@������������������������       �      ��       0����/#@������������������������       �               0#0# @�       �                   p��?/���?G       ";f�Q[@�       �                 h�/c?8&�_��?9       ]2� �U@�       �                 0VҼ?��צ��?       ��,[ufE@�       �                 @?�t:��?�?       m2 ��?2@�       �                    �?�KA<);�?       -mt��,@�       �                 P�T�?
�J���?       a���@�       �                 `	x�?�zœ���?       IG���t@������������������������       �               0#0#�?������������������������       �               z�5��@������������������������       �               0#0# @������������������������       �               ��#�� @������������������������       �      �<       ��/���@�       �                 �M��?��N3{��?       ]�9�+�8@�       �                    �?0&��:��?       ��0kk�4@������������������������       �               ��/���@�       �                 �fP�?�ѿ�FB�?	       G���W�)@������������������������       �               0#0#@�       �                  `s�?�`���6�?       /u��֝!@�       �                  ��??�@G���?       hu��@�       �                 pg��?|��`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @������������������������       �               0����/@������������������������       �               ��#���?������������������������       �               0#0#@�       �                 �Q�?�~���9�?       �q�Ί#F@������������������������       �               ��)��)C@�       �                    �?|��`p��?       �����@������������������������       �               H�4H�4@�       �                 ���?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?������������������������       �      ȼ       #0#06@�t�bh�hhK ��h��R�(KK�KK��h �B�  ���>��e@M��+c@���~�gb@�>��d@p>�c�^@L�dJ��P@�>��d@�����]@��+��+4@�>��d@M!Д[@��)��)3@�#����U@�-����@@0#0#�?��#�� @��On�(@        ��#�� @��On�(@        ��#���?��On�(@        ��#���?0����/#@        ��#���?��/����?        ��#���?                        ��/����?                D�JԮD!@                �cp>@        ��#���?                z�5��@                ��#�� @                ��#��@                �b:���S@鰑5@0#0#�?$�}��O@D�JԮD!@        Ip�}>@��/����?        ��#��@��/����?        ��#�� @                ��#�� @��/����?        ��#�� @                        ��/����?        �#���9@                ��#��@@��/���@        ��#��@@�cp>@                �cp>@        ��#��@@�cp>@        \Lg1��6@�cp>@        \Lg1��&@�cp>@        z�5��@�cp>@        ��#���?�cp>@                �cp>@        ��#���?                ;��,��@                ;��,��@                \Lg1��&@                <��,��$@                        ��/����?        ��#��0@��On�(@0#0#�?|�5��(@�cp>@        |�5��(@��/����?        z�5��@��/����?                ��/����?        z�5��@                �k(��"@                        ��/����?        ��#��@0����/#@0#0#�?        0����/#@0#0#�?                0#0#�?        0����/#@        ��#��@                �YLg1R@4����/S@vb'vb'2@��,���A@4����-O@#0#0&@�k(��2@��On�H@0#0# @��#�� @h
��F@0#0#�?        ���-��*@        ��#�� @��/���>@0#0#�?��#���?                ���>��@��/���>@0#0#�?;��,��@���-��@        z�5��@���-��@                ���-��@                ��/����?                0����/@        z�5��@                ��#�� @                ��#�� @�e�_��7@0#0#�?        �cp>7@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        h
��6@        ��#�� @��/����?                ��/����?        ��#�� @                ;��,��$@�cp>@0#0#�?<��,��$@��/���@        ;��,��@                ;��,��@��/���@        z�5��@                ��#�� @��/���@                ��/���@        ��#�� @                ��#���?                ��#���?                        ��/����?0#0#�?                0#0#�?        ��/����?        ��#��0@��On�(@vb'vb'"@��#�� @���-��@0#0#�?        ��/����?        ��#�� @0����/@0#0#�?��#�� @��/���@0#0#�?���>��@��/����?0#0#�?���>��@��/����?0#0#�?;��,��@        0#0#�?z�5��@                ��#�� @        0#0#�?                0#0#�?��#�� @                ��#�� @��/����?                ��/����?        ��#�� @                        ��/����?        ��#���?��/����?                ��/����?        ��#���?                        ��/����?        ��#�� @�cp>@0#0# @��#�� @��/���@0#0# @                �C=�C=@��#�� @��/���@0#0#�?��#�� @��/����?        ���>��@��/����?        ��#�� @��/����?        ��#�� @                        ��/����?        ;��,��@                ��#���?                        �cp>@0#0#�?        �cp>@                        0#0#�?        ��/����?        �k(��B@��|��,@�C=�C=@�YLg1B@0����/#@0#0#@��#�� @��/����?0#0#@��#�� @��/����?                ��/����?        ��#�� @                                0#0#@Ey�5A@��/���@        *�����;@��/���@        	�#���9@��/����?        ��#���?��/����?                ��/����?        ��#���?                z�5��8@                ��#���?                �,����7@                ��#�� @�cp>@                �cp>@        ��#�� @                z�5��@��/���@        ;��,��@                ��#���?��/���@                ��/����?        ��#���?��/����?        ��#���?                        ��/����?        ��#���?0����/@H�4H�4@        0����/@0#0#�?                0#0#�?        0����/@        ��#���?        0#0# @��#���?                                0#0# @        ��/���@0#0#�?        ��/����?0#0#�?        ��/����?                        0#0#�?        ���-��@                �cp>@;k�6k�G@        0����/@8k�6k�G@        ��/����?0#0# @        ��/����?                        0#0# @        �cp>@;�;�F@                k�6k�69@                0#0#�?                H�4H�48@        �cp>@��+��+4@        ��/����?                ��/����?��+��+4@        ��/����?0#0# @        ��/����?                        0#0# @        ��/����?vb'vb'2@                vb'vb'2@        ��/����?                ��/����?        z�5��(@��|��<@�6k�6�S@        0����/#@0#0# @        0����/#@                        0#0# @z�5��(@0����/3@��jS@z�5��(@0����/3@�+��+�K@z�5��(@E�JԮD1@��8��8*@\Lg1��&@��/���@H�4H�4@[Lg1��&@        H�4H�4@z�5��@        H�4H�4@z�5��@        0#0#�?                0#0#�?z�5��@                                0#0# @��#�� @                        ��/���@        ��#���?���-��*@��+��+$@��#���?���-��*@H�4H�4@        ��/���@        ��#���?�cp>@H�4H�4@                0#0#@��#���?�cp>@0#0# @        �cp>@0#0# @        ��/����?0#0# @        ��/����?                        0#0# @        0����/@        ��#���?                                0#0#@        ��/����?��-��-E@                ��)��)C@        ��/����?0#0#@                H�4H�4@        ��/����?0#0#�?        ��/����?                        0#0#�?                #0#06@�t�bubh,h-ubh8)��}�(h;h<h=h>h?Nh@KhAKhBG        hChShDNhEJ�%hFG        hGNhHG        hKhTKhUhhK ��h��R�(KK��h �C              �?       @�t�bh\hihlC       ���R�hqKhrhuKhhK ��h��R�(KK��hl�C       �t�bK��R�}�(h?KhK�h�hhK ��h��R�(KK녔h��Bh3         �                  ����?h^�TS�?,      @�g�}@       a                 @���?ZsԪt�?�       ����m]r@       :                 �l�}?�*��m��?n       �V�=%f@                        ���b? ��7 �?B       Wt���[@                         �3��?t;�cqW�?       e��"!A@                        @Ws�?:�c3���?       �uk��1@                            �?�O-r��?	       �.w��e)@������������������������       �               0����/#@	       
                 �ȊV?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ��#�� @������������������������       �      �<       ;��,��@                        `�Z?��i�@M�?       ���wzb0@������������������������       �               ���-��*@                         m�a?j%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?       -                 �G�s?�L�]�?0       �A�E#~R@       "                    �?�}Cl��?$       �(q��K@                        @��>(#����?       z�߄�C@������������������������       �               ��/����?                        `��?ԇQ_���?       �'3�	C@������������������������       �               z�5��(@       !                 `�ռ?l\Cl[��?       =�s�d�9@                        `�yU?�q���?       ��|�^1@                        �߯�> �=�Sο?
       ����,@                         Pmj�?�d�$���?       �T�f@������������������������       �               ��#��@������������������������       �      ȼ       ��/����?������������������������       �      ��       �k(��"@                          Џ~�?^%@�"�?       ��[�@������������������������       �      �<       ��/����?������������������������       �               ��#���?������������������������       �               ��#�� @#       $                 �/��?�����?       ��X�)B0@������������������������       �               ��/����?%       *                 �H/?X����?
       P	K��,@&       '                 ����?�����?       ��X�)B @������������������������       �               ;��,��@(       )                 _5?`%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?+       ,                 �7�?      �<       z�5��@������������������������       �               ��#���?������������������������       �               ;��,��@.       3                    �?���3�g�?       ص5��2@/       0                 �.�?\n����?       � ��w<@������������������������       �               ��/����?1       2                 жd|?�d�$���?       �T�f@������������������������       �               ��/����?������������������������       �               ��#��@4       5                 �m�?�L����?       Yk���>)@������������������������       �               ��#���?6       7                  y��?�F���?       :�.�-'@������������������������       �               ��/���@8       9                 �j%?Ĕfm���?       ��Z�N@������������������������       �               �cp>@������������������������       �               ��#���?;       X                 �6��?�|�)��?,       ����;Q@<       S                  �/�?�Skc���?$       �n�laM@=       P                 �Uu�?��o8��?       ��Z��H@>       I                  %�r?0�|�5�?       ����^E@?       F                 �.KR?��߭Q��?       �QVl�0@@       E                 `�J?��k*���?
       ���b-@A       D                 @F�`n����?       � ��w<@B       C                 ��=�?f%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               z�5��@������������������������       �      ��       E�JԮD!@G       H                   �P�?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?J       K                    �?8r�]i��?       ��U�i�9@������������������������       �        
       鰑5@L       M                 ny�v?( k�Lj�?       �q��l}@������������������������       �               �cp>@N       O                 PeT�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?Q       R                 p���?�AP�9��?       i��6��@������������������������       �               ��/����?������������������������       �               ��+��+@T       U                 �~(�?�K��t�?       L����"@������������������������       �               z�5��@V       W                 h��?v��`p��?       �����@������������������������       �               0#0#@������������������������       �      �<       ��/����?Y       `                 �/��?����?       ���"�X$@Z       _                 (/��?޺W�w��?       �'DQm"@[       \                 Ш��?��6L�n�?       �E#��h @������������������������       �               ;��,��@]       ^                 `�S?bn����?       � ��w<@������������������������       �               ��#�� @������������������������       �      �<       ��/����?������������������������       �               0#0#�?������������������������       �      ȼ       ��/����?b       �                 �7a?QUl_���?R       �F<+]@c       �                 ����?<3$���?;       �k-C�T@d       �                  �~��?�O�I	�?-       ��W���O@e       �                 �
h�?\������?       �r��E@f       q                 0�2�?vx�r��?       ���a��@@g       n                 ��Yk?B�%lX�?       ��f�B�-@h       m                  ��?����e��?       �ga��!@i       j                     �?d�r{��?       e�6� @������������������������       �               0����/@k       l                 �qʌ?b%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               0#0#�?o       p                 (I��?T����1�?       ��;9�@������������������������       �               0#0# @������������������������       �               ��#��@r       y                  �9��?�W�w��?       �'DQm2@s       v                 @2�?h�s�	�?       f���*@t       u                  pS��?      �<       \Lg1��&@������������������������       �               ��#��@������������������������       �               ���>��@w       x                 8<o�?���/��?       V��7��?������������������������       �               ��/����?������������������������       �               ��#���?z       }                 ��ȕ?П��X�?       m�n�/@{       |                 `U�?|��`p��?       �����@������������������������       �               0#0# @������������������������       �      �<       ��/����?~                           �?      �<       ��#�� @������������������������       �               ��#���?������������������������       �               ��#���?�       �                    �?d)���?       y��uk!@������������������������       �               ��#���?������������������������       �               ��/���@�       �                 p
E�?���~�w�?       X��]��5@������������������������       �               �k(��2@�       �                  4W�?���`p��?       �����@������������������������       �               ��/����?������������������������       �               0#0# @�       �                 @���?�Rn*l�?       6���2@�       �                 ��|�?P��W�?	       94���%@������������������������       �               ��#���?�       �                  ��d�?���k�L�?       sk��#@�       �                   ��?�LU���?       h�ҹ^�@������������������������       �               0����/@�       �                 �G��?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?�       �                 0釵?�J���?       ��*]Y @������������������������       �               0#0#�?������������������������       �               ��#���?������������������������       �               0#0# @�       �                  �p{?��Ɵ��?       �(�NA@�       �                 ���?d����?       �����!@�       �                 n�x?�v�;B��?       ՟���	 @������������������������       �               �C=�C=@������������������������       �      ȼ       ��/����?������������������������       �      ȼ       ��/����?�       �                 ��C�?�-�bƲ?       =�7*9@������������������������       �      ��       ��+��+4@�       �                 @��?�@����?       ���a�@������������������������       �               ��/����?������������������������       �               0#0#@�       �                 @�ޏ?�Cg�b*�?l       X"QQGf@�       �                 ��=�?�*A��$�?G       �����]@�       �                 H<��?�q=����?*       �A�錁P@�       �                 `�ۊ?z=:�BY�?       �J�C@�       �                 p��z?���5�?       D�)�B=@�       �                  ���?��<��?       v=�x�8@�       �                 ��Qg?�q���?       ��|�^1@������������������������       �      ��       {�5��(@�       �                 ���T?4=�%�?       �(J��@������������������������       �               �cp>@������������������������       �               ��#�� @�       �                 f�?      �<       ���-��@������������������������       �               ��/����?������������������������       �               �cp>@�       �                 (�s?      �<       ;��,��@������������������������       �               ��#���?������������������������       �               ��#��@�       �                 @�C�?nQ��?       �s�=�!@������������������������       �               ���-��@������������������������       �               ��#�� @�       �                 0�2�?n�4$�?       �,'{�;@�       �                   ���?f�q����?       O�Q*s�/@�       �                 ීv?�� ��?       rp� k@������������������������       �      �<       ��/����?������������������������       �               0#0#�?�       �                    �?�n���k�?       3��&�*@�       �                 ��z�?Hy��]0�?       ���y"@������������������������       �               ��/����?������������������������       �               ��+��+@������������������������       �               �C=�C=@�       �                 `��?�\U�?       �{����'@������������������������       �               ;��,��@�       �                 �Q��?��[����?       Hl�_A@������������������������       �               ��/���@�       �                 �p�?z��`p��?       �����@������������������������       �               0#0#�?�       �                 �$G�?|�G���?       ��%�|�?������������������������       �               0#0#�?������������������������       �      �<       ��/����?�       �                   p��?��2�6�?       %����J@�       �                  ���?�5�n ��?       ��/�@@�       �                 P�?n'1n 6�?       E��N:@�       �                 ����?��Dr�?       �9[�7�!@������������������������       �               0#0#@�       �                 �]!�?$ k�Lj�?       �q��l}@������������������������       �               ��/����?�       �                 ��ϣ?`%@�"�?       ��[�@������������������������       �               ��#���?������������������������       �      �<       ��/����?������������������������       �               S2%S2%1@�       �                    �?��r�g��?       ��1ֻ�@������������������������       �               �cp>@�       �                 ����?T����1�?       ��;9�@������������������������       �               0#0#�?������������������������       �               ��#�� @������������������������       �               ��-��-5@�       �                 X�*T?�TT2S�?%        n�K�M@�       �                 ��x�?fQ��?       �s�=�!@������������������������       �      ��       �cp>@�       �                  ���?\n����?       � ��w<@������������������������       �               ��#���?�       �                  P˗?���/��?       V��7��?������������������������       �               ��#���?������������������������       �      �<       ��/����?�       �                 @55�?�(.�?       Q��I@������������������������       �               H�4H�48@�       �                 ��t�?�N�+�?       ����:@�       �                 @f*�?�T`�[k�?	       �m����0@������������������������       �               ��/����?�       �                 �N��?��E�B��?       dߞKC.@�       �                 ��ݻ?�� ��?       rp� k@������������������������       �               ��/����?������������������������       �      �<       0#0#�?������������������������       �               H�4H�4(@������������������������       �               vb'vb'"@�t�b�Q      h�hhK ��h��R�(KK�KK��h �B  y�YLGc@鰑Nc@�N��Nld@��>���^@K!�M\@�s?�s?M@��k(/T@��]�ڕU@��+��+$@%�}��O@�'�xr�F@        �k(��"@��On�8@        ��#�� @0����/#@        z�5��@0����/#@                0����/#@        z�5��@                ��#���?                ��#�� @                ;��,��@                ��#���?��/���.@                ���-��*@        ��#���?��/����?        ��#���?                        ��/����?        ��b:��J@%jW�v%4@        �,����G@��/���@        ��,���A@��/���@                ��/����?        ��,���A@�cp>@        z�5��(@                [Lg1��6@�cp>@        ���>��,@�cp>@        ��b:��*@��/����?        ��#��@��/����?        ��#��@                        ��/����?        �k(��"@                ��#���?��/����?                ��/����?        ��#���?                ��#�� @                {�5��(@��/���@                ��/����?        z�5��(@��/����?        z�5��@��/����?        ;��,��@                ��#���?��/����?        ��#���?                        ��/����?        z�5��@                ��#���?                ;��,��@                z�5��@��On�(@        ��#��@��/����?                ��/����?        ��#��@��/����?                ��/����?        ��#��@                ��#�� @鰑%@        ��#���?                ��#���?鰑%@                ��/���@        ��#���?�cp>@                �cp>@        ��#���?                ��,���1@�)�B�D@��+��+$@<��,��$@������C@vb'vb'"@���>��@�+Q��B@��+��+@���>��@����z�A@        z�5��@鰑%@        ��#��@鰑%@        ��#��@��/����?        ��#���?��/����?        ��#���?                        ��/����?        z�5��@                        E�JԮD!@        ��#�� @                ��#���?                ��#���?                ��#���?��On�8@                鰑5@        ��#���?��/���@                �cp>@        ��#���?��/����?                ��/����?        ��#���?                        ��/����?��+��+@        ��/����?                        ��+��+@z�5��@��/����?0#0#@z�5��@                        ��/����?0#0#@                0#0#@        ��/����?        ���>��@��/����?0#0#�?���>��@��/����?0#0#�?���>��@��/����?        ;��,��@                ��#�� @��/����?        ��#�� @                        ��/����?                        0#0#�?        ��/����?        >��,��D@���-��:@J�4H�4H@=��,��D@�e�_��7@S2%S2%1@������C@E�JԮD1@�C=�C=@<��,��4@On��O0@��+��+@������3@E�JԮD!@��+��+@;��,��@���-��@H�4H�4@��#���?���-��@0#0#�?��#���?���-��@                0����/@        ��#���?��/����?        ��#���?                        ��/����?                        0#0#�?��#��@        0#0# @                0#0# @��#��@                ���>��,@��/����?0#0# @z�5��(@��/����?        \Lg1��&@                ��#��@                ���>��@                ��#���?��/����?                ��/����?        ��#���?                ��#�� @��/����?0#0# @        ��/����?0#0# @                0#0# @        ��/����?        ��#�� @                ��#���?                ��#���?                ��#���?��/���@        ��#���?                        ��/���@        �k(��2@��/����?0#0# @�k(��2@                        ��/����?0#0# @        ��/����?                        0#0# @��#�� @���-��@��+��+$@��#�� @���-��@0#0# @��#���?                ��#���?���-��@0#0# @        ���-��@0#0#�?        0����/@                ��/����?0#0#�?        ��/����?                        0#0#�?��#���?        0#0#�?                0#0#�?��#���?                                0#0# @        �cp>@=�C=�C?@        ��/����?�C=�C=@        ��/����?�C=�C=@                �C=�C=@        ��/����?                ��/����?                ��/����?H�4H�48@                ��+��+4@        ��/����?0#0#@        ��/����?                        0#0#@���b:@@�)�B�D@��8��8Z@Jp�}>@��/���>@�s?�s?M@��b:��:@�e�_��7@�A�A.@�k(���5@On��O0@        ������3@/����/#@        ���>��,@/����/#@        ���>��,@�cp>@        {�5��(@                ��#�� @�cp>@                �cp>@        ��#�� @                        ���-��@                ��/����?                �cp>@        ;��,��@                ��#���?                ��#��@                ��#�� @���-��@                ���-��@        ��#�� @                ;��,��@��/���@�A�A.@        �cp>@��8��8*@        ��/����?0#0#�?        ��/����?                        0#0#�?        ��/����?H�4H�4(@        ��/����?��+��+@        ��/����?                        ��+��+@                �C=�C=@;��,��@0����/@0#0# @;��,��@                        0����/@0#0# @        ��/���@                ��/����?0#0# @                0#0#�?        ��/����?0#0#�?                0#0#�?        ��/����?        z�5��@���-��@�
��
�E@z�5��@���-��@#0#06@��#���?��/���@��-��-5@��#���?��/���@0#0#@                0#0#@��#���?��/���@                ��/����?        ��#���?��/����?        ��#���?                        ��/����?                        S2%S2%1@��#�� @�cp>@0#0#�?        �cp>@        ��#�� @        0#0#�?                0#0#�?��#�� @                                ��-��-5@��#�� @鰑%@(S2%S2G@��#�� @���-��@                �cp>@        ��#�� @��/����?        ��#���?                ��#���?��/����?        ��#���?                        ��/����?                ��/���@'S2%S2G@                H�4H�48@        ��/���@#0#06@        ��/���@��8��8*@        ��/����?                ��/����?��8��8*@        ��/����?0#0#�?        ��/����?                        0#0#�?                H�4H�4(@                vb'vb'"@�t�bubh,h-ubeh,h-ub��e�memory�NhO�ub.