��c
     �imblearn.pipeline��Pipeline���)��}�(�steps�]�(�maxabsscaler��sklearn.preprocessing._data��MaxAbsScaler���)��}�(�copy���n_features_in_�K�n_samples_seen_�M��max_abs_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����f8�����R�(K�<�NNNJ����J����K t�b�C@     @V@      �?     ��@du��w@i�G5��7@�St$��@ffff&�@    ��@�t�b�scale_�hhK ��h��R�(KK��h �C@     @V@      �?     ��@du��w@i�G5��7@�St$��@ffff&�@    ��@�t�b�_sklearn_version��1.0.1�ub���gradientboostingclassifier��sklearn.ensemble._gb��GradientBoostingClassifier���)��}�(�n_estimators�K(�learning_rate�G?�      �loss��deviance��	criterion��friedman_mse��min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �	subsample�G?�      �max_features�N�	max_depth�K�min_impurity_decrease�G        �	ccp_alpha�G        �init�N�random_state�K*�alpha�G?������͌verbose�K �max_leaf_nodes�N�
warm_start���validation_fraction�G?��������n_iter_no_change�N�tol�G?6��C-hK�classes_�hhK ��h��R�(KK��h �C      �?       @      @�t�b�
_n_classes�K�
n_classes_�K�loss_��sklearn.ensemble._gb_losses��MultinomialDeviance���)��}��K�Ksb�max_features_�K�estimators_�hhK ��h��R�(KK(K��h�O8�����R�(K�|�NNNJ����J����K?t�b�]�(�sklearn.tree._classes��DecisionTreeRegressor���)��}�(h9h:�splitter��best�h@Kh;Kh<Kh=G        h?NhGNhD�numpy.random._pickle��__randomstate_ctor����MT19937���R�}�(�bit_generator�hr�state�}�(�key�hhK ��h��R�(KMp��h�u4�����R�(Kh!NNNJ����J����K t�b�B�	  C�&+�cCI�o��乾y_m?��Yf���"H�֝�2T��v�B��h��iC�˾��܃�5�!z��w�]�1�L�d�)�[6�r��Y�/������9tGxq-���K�#�_��_ 4},,������៩sz� �b�#��������5�����	z^����LA¨f�Et0kD-1�wK�����vB��ī)��Odر_�	�sA��X�'��iWH��yd�9�Gk�Wc��!o@pm�{�Z>тx ���e����=��A}>s�*e�-�J=D˼,���]�:6�]����YB@L�@(ΰ�+���5�%�&dE���'�ko��K��}?�h�#���ӕe�aB)5�=6__��c�d��}!ds�� �H厍�V�m�l2y�
��~#�ꤩ|��Vvcc	F��E6��]'iө!|<o�f�	֒��9�`ð𖼮
�O�Wf@�*�0���<K�$(�o�s�ǋ��osQmM���3�I9m��e�Z���	,oes"jE0���庺R����� ���C�X\�j�sX�WǍ9�I�`�Ū�7��fZ;�<�k1���g�Tb��Epnh(L��J3m�K��ů�;�U^,�]Ґ%�(ø�lw���#�O��=�.�Q	h�w��_���/�W�a�Ě�1y�b�b-������8g�@�2O�J�V�ïpg�(,4�UX���t���r�9{���Jز`9�G|���|{�-��G���M�����I��q���#EAl�o�5�d�[$#�4�C&=o!�wf}�J�J5���&�_�7H����k��)M�/���8^sV���#ZKDS";�[����P�s�" !���(:��AIq���IY ��������վ��l[��G��ܢ�]P��!;O�ԁ�ԛ衭��jJ�I��K��J�*k��c�X�;�i�i������-H�s�<D��)yX��x��V�b��	�e5�ڵ���v�����$�2�b��%!Fdj��)��5�>F@��b[�/NG)��YJ��֍�5A��4�  9�3C!�YO�5~��%�꛸�ƨ��i���ɩ.~�Mi�t���.(��傚0�c%��	�m�؁"H��� G�+[�6�ҙ�0g'xy_L���m7���gX�}���W'����o�;��nL�~�L�}5@��҄}#�D��"�j_�k�k�ޢ!������e�G��2�?>��㒠	����лg?�<�	�����(�l���__闸>�EQD�P��.��c�ո`�GUB��9�mg��Җ�#k+2�`K��O�S�ߺ��xz���]B�	�)x�)�CI�e���AiN����T~Mx���^T�c̜:���g�2DGVf�M���	)����c��*��|�vy{0E5��ΐ��0GaO_2�Է�27iQ���xb��!k� �p,��NR\d��}P%	�-��g�����c\�@6_�3��k��5Ї��~�(1�*�"Z�L�Gv��̹Q�*B3�CD�� }�|�p{��לZ��j�[�g�];�?�N;����ś q�\�@s�?q+��x�T�GӔU!�7/�_��h<�Q��!;;9�c�@�{R{�ˢ�(�ڵ�(�/>ւ��c�Jif�T@�\�7�j.��7t��w���"g����VeGA������y��;x|��y퀈7A����DA|)����qr�b���O ��棏ZeJ$����U<#��(]�ٍRo�1��#�|S���#�UWM��W�~�}��m���7Y�@{�d[h1(����V��^��Mq�%�B�z[~
��F3p�ȓm��?���ǖKy?�_"�Zc��ע �fh}��o��q�N��l+���^��wm��q��n�y;�_���h�? �nJ��A+u�U�`X��s�J�h�&sq���9}�W�/�'!����RJ�'`������ݼ^�Q3��@ɼ�(�tJP�� �h��°��-cKmiSfV���iz�.�Y�3��]r6?@P���]��ʆj�pM�]��|��:��>g�E4��W 9)aD3�0��Q�I1���^[P!�~uk�=��I�K�ɝ?:5l���)��Y"�	 ���.�Z�<?�~�)uu91#��޿&"`��1��v�������<���+�d�:6>î����6�a�����Z��8�mv��.)+����D�ܱC��6�cr�� �8%Fx�/�0B�[΂V�/0X6�4 V�}��<�((6!�E�ڈ�B����Z�cԏ�����t�S� )�jt��"M^/i���fe��-i5���<��O��W:��E����>J�q����E�qR<�7ie1���e�d����,���c'�_h DMþ�p�t�*�Q�F/��.Ҵ�!�8� B�\�uy��^�F7�[� �{���خ��[��4�uZqB���hÀ%E��$������=���vO���Z�M�k���q�h�n�	_U_B��t�b�pos�Kxu�	has_gauss�K �gauss�G        ubhAG        �class_weight�NhBG        hK�
n_outputs_�Kh\K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h�i8�����R�(Kh!NNNJ����J����K t�b�C       �t�bK��R�}�(h@K�
node_count�KK�nodes�hhK ��h��R�(KKK��h�V56�����R�(KheN(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(h�h�K ��h�h�K��h�h�K��h�h K��h�h K ��h�h�K(��h�h K0��uK8KKt�b�Bh         .                 P7&E?�e�,��?�           �}@       !                 @�Ц?�!I���?           �q@                        ����?	k��9�?�             l@                        �$?Z?�*;L�?x             ^@                        ��IL?�q�q�?             5@                        ����?�q�q�?	             "@������������������������       �      �?              @������������������������       �      ��             �?	       
                 �1?�8��8��?             (@������������������������       �      p<
             $@������������������������       ��������?              @                        P �s?GS%��?c            �X@                        �U���T%ޑ��?F            �Q@������������������������       �     �?             8@������������������������       ���nkK�?.             G@                        �i�?�f7�z�?             =@������������������������       ��	j*D�?             *@������������������������       �    ��?             0@                        p�%h?RN���?i            @Z@                        0�2�?!{��e�?5            �J@                         �\�?�����H�?-            �F@������������������������       �Y�<ݚ�?	             "@������������������������       �������?$             B@                         �t�?�������?              @������������������������       ��q�q�?             @������������������������       �      �<             @                             �	j*D�?4             J@                        `��?��G�z�?(             D@������������������������       ��q�q�?             @������������������������       ��t����?"             A@                            �?/�q�q�?             (@������������������������       �                     @������������������������       ��q�q�?             @"       )                 �H�9?d�� ż?>             O@#       (                  @���?��}b~|�?9            �L@$       '                 @���?N4և���?8             L@%       &                    �?�1�`jg�?7            �K@������������������������       �q�q��?             2@������������������������       �      �<%            �B@������������������������       �     ��<             �?������������������������       �      ټ             �?*       +                 `�C?���Q��?             @������������������������       �                      @,       -                  ���?�q�q�?             @������������������������       �                     �?������������������������       �      p<              @/       B                 `9�`?�?�C+�?�             g@0       =                 ��U�?�'݊U�?C            �P@1       6                  �/�?�����?&             C@2       5                 `�Z?~X�<ݪ?             2@3       4                  Џ~�?      �?              @������������������������       �                     �?������������������������       �      �<             �?������������������������       �      p<             0@7       :                 ��D�?�G�z��?             4@8       9                 �_�j?�z�G��?
             $@������������������������       �      �?             @������������������������       �      �<             @;       <                  �E�?��G�z�?
             $@������������������������       ������H�?	             "@������������������������       �      ��             �?>       ?                 �|�?JB���?             =@������������������������       �                     :@@       A                 H�z�?�q�q�?             @������������������������       �                     �?������������������������       �      p<              @C       D                  ��~�?�w5�?v            �]@������������������������       �                     �?E       J                 p"�?      �<u            @]@F       G                 ��Ē?     ��<d             Y@������������������������       �      �<1            �H@H       I                 p��?     ��<3            �I@������������������������       �      �<1            �H@������������������������       �     ��<              @������������������������       �     �ݼ             1@�t�b�values�hhK ��h��R�(KKKKK��h �BX  �<�"h8y�O%x��S�?51��^�?�%�2��?��F($�?K�O�v�?��F���?wwwwww��x��οxwwwww�;V ��c�?hi�i��?V K����?�I���?�����??(��5��?�fy{�k��d�/X��?�W��,�?k� O��0Y}���ʿ�~�	��?�'���쿠���c�?�1^��?��#�� @���ڐ��?��!���?�1^��?Eٰ`�?��F($�?wwwwww�e���a��?;,tG�ȿ�T�Ϳ;����	п�Z�هѿ�e4��\޿ywwwww���#�� @��#�� @HU2��?��#�� @��F($�?��#�� @wwwwww�ɡ����Ͽ���ob��Y�v���y�|��-�ѿA�Iݗ��?��#�� @wwwwww�wwwwww￦)�C�-�?��~������F���?wwwwww���!���?�<����?wwwwww���7�<gҿwwwwww���F($�?��#�� @wwwwww�u_[Կ��#�� @V[4�ԿO[4�Կwwwwww�^[4�Կwwwwww�wwwwww�wwwwwwￔt�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KEh�hhK ��h��R�(KKE��h��B         2                 �6Sz?�&��?�           �}@                        ��??k���X"�?           �w@       
                 @�W?4�X���?           �p@       	                 ��IL?���!pc�?             6@                        Pu�?�eP*L��?             &@                         ���?�q�q�?	             "@������������������������       ��q�q�?             @������������������������       �q�q��?             @������������������������       �                      @������������������������       �      ��             &@                          �G�?�&z�,�?�            @n@                        �С?џ[;U��?             =@                        ��GA?\X��t�?             7@������������������������       �                     @������������������������       �Y�<ݚ�?             2@������������������������       �      ��             @                        P��?Hb�3]�?�            �j@                        �v@�?��v>��?�            �g@������������������������       ��zœ���?�            `c@������������������������       ��eP*L��?!            �@@                        К��?�P�sײ?             9@������������������������       ��q�q�?             @������������������������       �      ��             6@       %                  �g<�?����� �?w            �]@                         �$I�?0�0�!��?3            �I@                         ��~�?X˹�m��?&             C@                        0�?      �?              @������������������������       �                     �?������������������������       �      ��             �?                         �X?X�<ݪ?$             B@������������������������       ��q�q�?             @������������������������       �pa�	�?!            �@@!       "                   ��?��
ц��?             *@������������������������       �                     @#       $                    �?�<ݚ�?	             "@������������������������       ��q�q�?             @������������������������       �                     @&       -                   p��?����� �?D             Q@'       *                  ����?C7�J��?7            �K@(       )                 ��J�?%��m��?             :@������������������������       ����|���?             &@������������������������       ��r����?             .@+       ,                 �5P?����"�?             =@������������������������       �z�G�z�?             @������������������������       ��q�q�?             8@.       1                 �̑�?%�q-�?             *@/       0                  ��g�?      �?              @������������������������       �                     �?������������������������       �      ��             �?������������������������       �      p�             &@3       @                  �E�?:q�/��?Y            @V@4       9                  ����?���}<S�?.             G@5       6                 �%��?<a�	�?!            �@@������������������������       �      ��             >@7       8                 @���?#�q�q�?             @������������������������       �                     �?������������������������       �      ��              @:       ?                 �0J�?�θ�?             *@;       <                 �Th�?      �?             @������������������������       �                      @=       >                 �/�?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �      p<             @A       B                 �@�?      �<+            �E@������������������������       �      ��             8@C       D                 0�?      �<             3@������������������������       �      p�             &@������������������������       �      ��              @�t�bh�hhK ��h��R�(KKEKK��h �B(        ��^65����?s�M��z��l��N�?<��j�?k��2팿�<B��?�]�ῴ�/����?��/����?
�[,V��G�ͯg%�?�>��Z�?�bAs�X��e���?��/����?\�=���]k!>c����J�@ӿxS'6��?�b�ѿ�<B��?�bAs�X�F�v���?��f��w�?��)��Z�?��c+���?��/����?�bAs�X����?�<B��?�ArdF�?�P��r�?�bAs�X�jy�]��?Ft#uC����/����?A1�mv�?Ŋ��\�?;��&t\U�A�4�.�?�ė�%�	|-0�|�?v�DN��ۿP�N�B��?D�a%pPѿ��c+���?��/����?�bAs�X�bAs�X�֩��b\ӿ�Q��пXF�BLԿ�bAs�X�k��2팿��/����?�bAs�X��$nJ߽���c+���?�bAs�X���A��?�bAs�X��/����?�bAs�X�N�<ֿ�bAs�X�N�<ֿ�bAs�X�bAs�X�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KEh�hhK ��h��R�(KKE��h��B         ,                 ��g?h�;K�R�?�           �}@                        ��^�?'��v4v�?j           �v@                        0-3�?����W�?-           �r@                        (/��?�ְ�*�?�            `g@                        ��=�?�M��ȅ?�            @g@                        ��?p�W��#v?�             g@������������������������       �      �<�             f@������������������������       �����X�?             @	       
                 �/��?     �?              @������������������������       �                     �?������������������������       �      �<             �?������������������������       �     ��             �?                        �n�?A�q��?r            �\@                        0=�?�eP*L��?             6@                        @�Ap?      �?              @������������������������       �      �?              @������������������������       �      p�             @                         ��d�?V�Cc�?             ,@������������������������       ��q�q�?             @������������������������       �      �?              @                        �{��?�ܸb���?\             W@                          Y��?&-�_ .�?J            �R@������������������������       � �,���?C            �P@������������������������       �����X�?             @                         Z��?�E��ӭ�?             2@������������������������       �      �?              @������������������������       � ףp=
�?
             $@       '                 `'v�?Vu���?=            �N@       "                  �~��?��P���?)            �D@                           �?V�<ݚ�?	             "@������������������������       �                     @        !                 �؉�?y�G�z�?             @������������������������       �                     �?������������������������       �                     @#       &                  @���?0     �?              @@$       %                 ����?��a�n`�?             ?@������������������������       �                     �?������������������������       ���S�ۯ?             >@������������������������       �     ��<             �?(       +                 �00�?�������?             4@)       *                  pjS�?     �?             0@������������������������       �      �<             .@������������������������       �      �<             �?������������������������       �      ¼             @-       8                 �6Sz?��Q|ӭ�?n            �[@.       1                    �?և���X�?             5@/       0                 @M^i?�������?              @������������������������       �                     �?������������������������       �      ��             @2       7                 p�r�?�n_Y�K�?             *@3       6                 �Y�n?���!pc�?             &@4       5                 ����?     �?             @������������������������       �                     @������������������������       �      �<             �?������������������������       �      �<             @������������������������       �      Ƽ              @9       D                  �E�?�o�/��?Y            @V@:       ?                  ����?���}<S�?.             G@;       <                 �%��?�a�	�?!            �@@������������������������       �      �<             >@=       >                  `���?�q�q�?             @������������������������       �                      @������������������������       �      ��             �?@       C                 �0J�?��θ�?             *@A       B                    �?      �?             @������������������������       �                      @������������������������       �     �?             @������������������������       �      �<             @������������������������       �      ݼ+            �E@�t�bh�hhK ��h��R�(KKEKK��h �B(  'u_[��l���uqſn�y��yп���4 Կ�T��vԿ����Կg��Ao���A����pR���?0#0# @e��Ao��0#0# @�9X���Ŀ�Uv4���?0��Nʿ-T�LW�?f��Ao�￰��D���?gT�/n�?-�l?�?cL�V��Ϳ=���m�ѿ�W����"o}rXF��2Y}�����-T�LW�?���I9��ɪ�?Wj�v��?�k`�*�?e��Ao�ￛk�.&�?e��Ao��0#0# @2��}yl�?9HL�S�?e��Ao����,M�?e��Ao��`[4�����V'ѿf��Ao��0#0# @0#0# @tHRAT��?w@x��?4��}yl�?e��Ao��0#0# @6�泫?��h���h8�����?0#0# @e��Ao��e��Ao��0#0# @%�xK��?8�r ��?=�Pn;t�?3#0# @�S����?0#0# @e��Ao��L��?�pR���?0#0# @q�EϿ0#0# @0#0# @�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KGh�hhK ��h��R�(KKG��h��B�         2                  ���?�lj��?�           �}@                        ��a,?ǵ|��?4           @s@       
                  `���?�������?�            �c@       	                 ,&k�?<Q~� ǳ?             @                        ��h*?�/���?             @������������������������       �                     �?                        �h?�3�G�?             @������������������������       ���-��=o?              @������������������������       �0��"E�|?             @������������������������       �      p<             �?                         �P��?��I�z�?�            �b@                        Phd?`�'M��?C            �P@                        P]ڒ?'U/���?,             F@������������������������       �`+��O�?"             A@������������������������       �)<x�a�?
             $@                        T�@?J�L��Ω?             7@������������������������       �                     �?������������������������       �l���۞?             6@                          \��?���g��?T             U@                        \O̙?���љB�?             @������������������������       �                      @������������������������       �,�,:��?             @                        ��=�?�yU���?O            �S@������������������������       �W��qݡ�?             (@������������������������       ���8���?C            �P@       %                 P��1?
c�~��?�            �b@                         0?lg���]�?             @                        ��u?|�dF�?             @������������������������       �                     �?                        0z�?Ⱦ�6�p?              @������������������������       �                     �?������������������������       �      ��             �?!       $                  s��?薷����?             @"       #                 �j�? p/�u�>?              @������������������������       �                     �?������������������������       �      �<             �?������������������������       �      ��             �?&       +                 _5?��hK���?�             b@'       (                 h(�>?��@�t�u?             @������������������������       �                      @)       *                 ��K�? &G�M�D?             @������������������������       �                     �?������������������������       � h�Tp�?              @,       /                 P+�Q?�N�fs�?�            `a@-       .                 0�̇?|�3t^�?             @������������������������       ���F1sW?              @������������������������       �      ��             �?0       1                 �l�e?�K��:"�?�             a@������������������������       �j�!�3��?             .@������������������������       ��|@b��?y            @^@3       4                 0��?�������?�            �d@������������������������       �                     �?5       :                 ���>*��g�ڤ?�            `d@6       7                  ���?(� A�t?             @������������������������       �                     �?8       9                 ����?�gj(�(T?              @������������������������       �                     �?������������������������       �      `<             �?;       @                 `��?I:<��j�?�             d@<       =                 �7�a?�"�����?             @������������������������       �                      @>       ?                  `<��?
� ��?             @������������������������       �`���J{?              @������������������������       �                     �?A       D                 �]t?��O��\�?�            `c@B       C                 �:?�}�*,�?             5@������������������������       �!��-Y�?             3@������������������������       �@$g���?              @E       F                  �z?��1#�?�            �`@������������������������       �ZQ�HG\�?	             "@������������������������       �Z�7�͖?}            @_@�t�bh�hhK ��h��R�(KKGKK��h �B8   �u$'Ϗ�Z�h�I?Г�D��?�7΃kƿa/^��xп��,CM��?�3-�p
տ���������ߋ����W��J�?i�����?�|���a�?�-�)��?�޵J���?�~��ސ�?�t�y�K~?�Ik�� ��<��*{�?�"�}3`e?ZPt��ֿ�Ik�� �W�=���@w���?FX���?�01i��e0'nY�����2/տ �៣y����,CM��?�b����ȿ�qoҁ�qA�HN��cשY�⿒����*�g��,��6����w�o\�}�wA�[���1�,��?C����?��d,�y�?���?�� ���?�������Ϡ.�ѿ����9�URR :��D�G�(����]5�n�?��y���ҿ	P�k;���q�v,N���ve������g���?a+���K�?"*R�X�?H`�#//�?C����?�Y�0+]��rB�ֿ�Ik�� ��'�����(����Z+}���P@�����-�q�?�)-�ѿ�?�(������O ���m ��R��i�ȵ�ܿ�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KQh�hhK ��h��R�(KKQ��h��B�         >                  �v�?��0,˴?�           �}@                        �jx?�o�\瞹?�            `l@                        ��v�?��_�;�?�             d@                        p�t?��h0���?�            `a@                        0���?8�iA�+�?�            �`@                        �U��?V��qĸ?x             ^@������������������������       ��7D���?o            �[@������������������������       �PZ0O�?	             "@	       
                 �,Ip?
}P
 :�?             ,@������������������������       � ��qԛ?             &@������������������������       �����h|�?             @                        pTF�?־�W|�?             @                         7�?.;�f�?              @������������������������       �                     �?������������������������       �                     �?                        ����?�����?             @������������������������       �  �C��z>              @������������������������       �      �<             �?                        ��9�?����-��?             6@                         H��? �/����?             @������������������������       �                     �?                        ���w?��Ա��?             @������������������������       �                      @������������������������       � �~1O�n?             @                        �i�N?nS���?             0@                        ���?h��.e i?             @������������������������       �                     �?������������������������       �                      @                        �c�w?���܍�?             *@������������������������       ���e�쀢?             @������������������������       ������W�?             @        /                 PFe�?n֏����?B            �P@!       (                 0�?�$��?3            �I@"       %                 P���?�,Z�[�?             6@#       $                 pD	�?ԫP��?             0@������������������������       �,[���?	             "@������������������������       ���-�ƨ�?             @&       '                 ��K?�F���?             @������������������������       ��O��n ?              @������������������������       ��7*�n5�?             @)       ,                 �5W�?\�Ĩ?             =@*       +                 X�)�?V4^J���?             @������������������������       �@۫�+q?              @������������������������       �      ��             �?-       .                 0Y�?f1;�ќ?             :@������������������������       �0ssu!��?             6@������������������������       �p�UO��?             @0       7                 �!�@?�n��^��?             .@1       4                 �ᒤ?�.��jf�?             @2       3                 0��?��yZ�u?              @������������������������       �                     �?������������������������       �      ��             �?5       6                 P'��?�t�����?             @������������������������       � �����`?             @������������������������       �                     �?8       ;                 �㨤?7���ǲ{?	             "@9       :                 ���?�/U�jzF?             @������������������������       �����oK?              @������������������������       �       �              @<       =                 @W�?�3��'?             @������������������������       ��Jp�һR?              @������������������������       �                     @?       @                 �$I�?�=���?�            �n@������������������������       �                     �?A       J                 ���?��.���?�            �n@B       I                 ���?3%B�p�?�             n@C       F                 q� ?�}Mub�?�            �m@D       E                   E(�?�3�d�Y�?             @������������������������       �                     �?������������������������       ��A�uVp?             @G       H                 pt"?e��$�?�             m@������������������������       �                     �?������������������������       �7$=G>�?�             m@������������������������       �     =             �?K       L                 pH�?n>E�!��?             @������������������������       �                     �?M       P                 �h�?6��t��?             @N       O                 ��^?����Sa?              @������������������������       �                     �?������������������������       �                     �?������������������������       �      8<             �?�t�bh�hhK ��h��R�(KKQKK��h �B�  $��b���?s-{k��?~$ҍ8w�?�C ;~�?��L�|�?R�Cw8t�?��OyB�?�
��̐�?I��!����S@�Ma���D}Kgx�?�ֈ}���?	9�R��?{�`މ2�n=���|�?){1�XK�?��`�Fx@����m�?�#]CZ��?�1PG9�?,��+��?��IeF9�?�'��@����?�W/A��?0N�К���;;)�4뿁�3�7�����o?�?��n��|�?;u�i7�?��f�s5�?h��I'(���/>S�����ԍ�ÿ��g�B�쿞ȁ@���kM��)��?��;���M������?V��sГ?+Cg���?�RM�&��?�c�[����Y������տ���*��?	�*���?�%��o�?%��-d�?LD��,�?A3HE;@��F��?&��t��?l��+���?���fƒ�X�a�6���1zĬ�翘c�[� ����}�?#�B��翐}=��?��+=⓿XG��?���'1���y�nS���6g<��i�M^;cɿ��`��
�>���?���`�Ho���j���?w�Y�+��C�I��nAsoc!ӿ����� ��Ӣ܇�ſ,w4��Ϳ?드17�*���k��c�[濔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KUh�hhK ��h��R�(KKU��h��B�         .                 ��\�?�Xq��R�?�           �}@                        �I�f?g�ː?5�?           �p@                        0�ǟ?w'���?�             n@                        ��9�?��?�v�?�            �j@                        �U����f�NP}[?�            �a@                        �R$X?`E̒O�R?8             L@������������������������       �P ���'.?             0@������������������������       � �k	P?(             D@	       
                  Y�i?���Z%]?W            �U@������������������������       ��wU�^>?:             M@������������������������       ��ƝƯm?             =@                        �Q�?uY��}�?F            �Q@������������������������       �                     �?                        �\ͥ?b)'��Y�?E            @Q@������������������������       ��8�|4�?             @������������������������       ��v	U�9�?B            �P@                        �m��?�j7��γ?             <@                        @?,�?��˼��?             @������������������������       �                     �?                          E(�?4��qJ��?             @������������������������       ��/��=�?             @������������������������       ���/O��?             @                        `f�|?(����?             5@                        @b#�?��>t}�?              @������������������������       �                     �?������������������������       �      �<             �?                        �a��?�
�q�?             3@������������������������       ��An{�>f?             2@������������������������       �      �<             �?       +                  <��?�ةyYs?             :@       $                   ��?��{~�l?             8@        #                 pW�~?Ue@��;s?             @!       "                 �@�? i^����>             @������������������������       �                     �?������������������������       � \�B2�>              @������������������������       �      @�             @%       (                 ��;�?���gHa?             2@&       '                 �h�? J�*'�1?             .@������������������������       � ��ĭ�>             ,@������������������������       �      ��             �?)       *                 b4�?G��&�~?             @������������������������       �                     �?������������������������       �      @<              @,       -                 Nq��?��i�GB?              @������������������������       �                     �?������������������������       �                     �?/       8                   \��?�4N�K�?�            �i@0       7                 �0H�?��Aj��?(             D@1       6                 (;�?0�-�ԁ?'            �C@2       5                 0n1�?hNSw|?#            �A@3       4                 �^<:?d���av?!            �@@������������������������       �H�ކ[�?             2@������������������������       � r�u97?             .@������������������������       �      p�              @������������������������       �                     @������������������������       �      ��             �?9       H                 �{��?����o�?�            �d@:       A                  ;�?��pH�?F            �Q@;       >                 �!�?w{J�W�?             @<       =                 P�ټ?	_�'{w?              @������������������������       �                     �?������������������������       �      0�             �??       @                 p[R�? ��ubC?              @������������������������       �                     �?������������������������       �      �<             �?B       E                 `Fe�?��)����?B            �P@C       D                 �\3�?JV>	^g�?5            �J@������������������������       �z�nu��?             3@������������������������       �R�����?"             A@F       G                 ���?XȦ���?             *@������������������������       �������?             @������������������������       �h&��bf?
             $@I       P                 �\��?I_�UQ�?_            �W@J       M                 Ш��?M�J&!�?Z            �V@K       L                 �0Mt?"�\ZG��?             *@������������������������       �h]"�?              @������������������������       �      P�             @N       O                 �Ϻ�?�Mr�l��?M            @S@������������������������       ��v�J`�?              @������������������������       �r_�>�?K            �R@Q       R                 vX�_?]Ɨ��l�?             @������������������������       �                     �?S       T                 V�"�?`���Q݂?             @������������������������       �                     @������������������������       �      p�             �?�t�bh�hhK ��h��R�(KKUKK��h �B�  0Ӯ����!�e�l��Ƥ��ɳ�Ձ}#ڑ���{=ۤ���F_�춿��������P[����������L���BP �~���ێk�����-�N���%�ܼ8޻��ăF&!�?�HSmX�{J�^�u?j���4�?��U���!@���?5�"�ӈ���m��?�P���EXh��?E���e�?	����?,�w!ɐ��t_��:迪�娐b�f�)�N��?��@u�?L�r}��?$�R�{�����y��@��7X�
6GK#q�?�i��䙵? ��<^v�?.��a8|�?ߚ���:�?�ƍ.�?ִ��6GK#q�?�|y&j�����y���z6]��-���B�?b�A����\z�T���"����T��E�O�����Ѐ�	�Y7���
6GK#q�?	6GK#q�?.��t&6@�6H�/��?�a\����?bC�x@~�?X�_�'�?
6GK#q�?�zY!��h�W��	�?[����@|��w��@M����?U3��?�O��u��?��e��n�?�M����?��^f�?y�|��?�~��+�?o��7�?��K鼿�;M����6GK#q�?����Nh�?�>�_q��?Ꜵ�`�?"-��!��?/�Τ5S@��5��?6GK#q�?��оP��?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KSh�hhK ��h��R�(KKS��h��B(         :                  �=�?a��J(�?�           �}@                        p۶�?��j��?            q@                         �ڦ?_�Q��b�?�            �k@                        @&ɥ?
."����?�            �b@                        ����?OTWǢ?�            @a@                        ��??��,6�J�?            �_@������������������������       �λM΋�?^            �W@������������������������       �v�,�):�?!            �@@	       
                 �4�r?�b8�h�?             &@������������������������       ��j"$G�?             @������������������������       �7L2r�R�?             @                         �J�?N<�G�?             &@                        ����?b?Gfd�?
             $@������������������������       �<
^$ju?              @������������������������       � N�@�q?              @������������������������       �      ��             �?                        ��Yk?��$0���?I            @R@                          ҏ�?Ys�Pjf�?!            �@@                        �j5?�j҂n�?             @������������������������       �B�]NU�?              @������������������������       �     �`�             �?                         �\�?>�a�]�?             >@������������������������       ������ū?              @������������������������       ��Ż=N&x?             <@                        ����?�-!)�?(             D@                        �$�?����?"             A@������������������������       �s7c9���?             4@������������������������       �F��I'-W?             ,@                        ���?$�:3�m�?             @������������������������       ��vM�|e?             @������������������������       �xY���>              @        -                   s��?K�A�5�?4             J@!       &                 xv�Q?�����Ŕ?             :@"       #                 K)w?�v����?             @������������������������       �                     �?$       %                  I<�?8��S��?             @������������������������       �����g?              @������������������������       �      T<             �?'       *                 �lO�?�Y�q���?             6@(       )                 ���?�	�_[p?             (@������������������������       �p�Z��h?             &@������������������������       �     p��             �?+       ,                 ��?������?
             $@������������������������       �:��ј�?	             "@������������������������       �                     �?.       3                  �^�?�i�]�?             :@/       2                  As�?0��e��?              @0       1                 �}��?�֢��w?             @������������������������       �j�[�e�m?             @������������������������       �����V?             @������������������������       �      p�             �?4       7                 �p�?��P�)5�?             2@5       6                 h��1?�&+���?             @������������������������       ����	f2T?              @������������������������       �                     �?8       9                 p��?XM�r�\z?             .@������������������������       ��D�v�l?             ,@������������������������       �     �<             �?;       R                  @���?U ��2��?�            �h@<       C                 ��ځ?��TY{�?�            �h@=       B                 �5�z?E����?             @>       ?                 P��?�o�hb�?             @������������������������       �                     �?@       A                 l�Y`?@�`+X�6?              @������������������������       �                     �?������������������������       �       �             �?������������������������       �      �<             �?D       K                 `��?�S�+ˈ?�             h@E       H                 �ڡ3?�ϵ�i�?             *@F       G                  v�?��=5ݔ?             @������������������������       ��s��&3r?             @������������������������       �F�*�C�[?              @I       J                 ���{?�8�"PC?              @������������������������       �                     �?������������������������       �X��Hĭ?             @L       O                 ����?����CG�?�            �f@M       N                   �P�?zP1��?�            �a@������������������������       ��a�?� �?2             I@������������������������       �*xЇ��|?[            �V@P       Q                 ЩI�?�C�M	h?'            �C@������������������������       �                     �?������������������������       �U��4�`?&             C@������������������������       �     ��<             �?�t�bh�hhK ��h��R�(KKSKK��h �B�  ��`vt?�|���ѝ?�oxXo�?��譡?��[�Uޔ?׌˭�c�?Z$���?z�e�ۿ�kt)���4��=:�?�,��������$�?P�\S�6�?<ҞE���?X�Zd�o�?��x�Lz�?RT>�Ht��I0���Y��kZп�߄���4�����忑��Ǚ����F�?v�HB�5��+��ؐ?.��S]{�*�g�3�?�z<`1��)�����?��SW��?��B=��V��r���?��R$l�?e@'\*�ĿX���?��{��o;����[��H����L��?��xh1:�?�,�񁇹?=j���%�?��)e'��>�uBvB�?�CG]��?v�2a�J�?�`4�0��?���c��?^:�!^�?c�:�t�?�zd���?�����鿲o����?��rC{��?KUŨ��?�Զv�@�$�z��?���K�:�?�����;������#[}�����	ſ��U��p�?�$*�?.�G%ˬ�y�!:��񆶞#+��-Ha�0�ma������^���ڹ���PN�˿�������CD�[�H՜�p��)��nf�i��.��忆�oU�����T���6�񹒲?;�|��׿~~%�_ѧ�e��N��Z�G��z翳�7$���?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KSh�hhK ��h��R�(KKS��h��B(                            �G�?��"n�?�           �}@                       ��z�?:{�}&Y�?@             P@������������������������       �                     �?                        ���u?� �d-�??            �O@       
                   ҏ�?(Zm��|�?             5@       	                 �.s�?@X��ؙ?             4@                        ��H�?d���ͳ�?             3@������������������������       �o��11�?             .@������������������������       ���ү��?             @������������������������       �      ��             �?������������������������       �      ��             �?                         ?Dy?H������?*             E@                        �;�?�~�M���?             @                        ����?��[�c?              @������������������������       �                     �?������������������������       �      `�             �?������������������������       �      ��             �?                        ,*���x)T���?'            �C@                        ��0�?�{j��ё?             (@������������������������       �����
Ď?             @������������������������       ���KW}?             @                        �$I�?3��?             ;@������������������������       ���x�>�?             4@������������������������       ���h2�g?             @       6                 ��n�?���4�x�?�           �y@       )                 p۶�?5_8
�.�?�            `o@       "                  �Mm�?y�	P�d�?�            `i@                         ���?w��4�?�            �e@                         �P��? �jњ�?�            �c@������������������������       �[���XD�?,             F@������������������������       ���\.�?q            @\@        !                  �J�?.����?             2@������������������������       ����(�r?             1@������������������������       �      �<             �?#       &                 P�bf?�8����?             <@$       %                 ��l?��{�9��?             .@������������������������       ��#A_�ō?             @������������������������       ���.���?	             "@'       (                 �)p�?����b?             *@������������������������       ��|1�)x6?              @������������������������       ����aUP?             &@*       /                 �-�?>�����?0             H@+       .                    �?T���y�?             @,       -                 �R�?��gj�4f?             @������������������������       �������?              @������������������������       �      `<             �?������������������������       �                     �?0       3                  �^�?,���^�?,             F@1       2                  As�?ӫ~86܂?             ,@������������������������       �W�-PȀt?             *@������������������������       �      �<             �?4       5                 p��?���mwv?             >@������������������������       ���t��p?             7@������������������������       �p����j?             @7       D                 ���?FZ��i�?�            �c@8       ?                 �
�?ZJΧ��?             (@9       <                  �Q�?g �1�ǡ?	             "@:       ;                 ����? � �?              @������������������������       �                     �?������������������������       �      h�             �?=       >                 �>�?��;�ļ�?             @������������������������       ��Ud7Y��?             @������������������������       �$o�׼X?              @@       C                 t��A?И��̮?             @A       B                �o|?@kQ��Ґ?              @������������������������       �                     �?������������������������       �      �<             �?������������������������       �      ��             �?E       L                 pZ9�?�?4Ğ?�             b@F       I                 �O�??����?1            �H@G       H                  �P�?��XdӼ�?
             $@������������������������       �                     �?������������������������       �(ؐ�o?	             "@J       K                  �u��?$�2��?'            �C@������������������������       �IL$��?%            �B@������������������������       ���C�[6�?              @M       P                  ���?�,��O��?`             X@N       O                 ��\�?0cXJ�,�?              @������������������������       �                     �?������������������������       �      �<             �?Q       R                  �@�?�ȓd��?^            �W@������������������������       �{�j���?]            @W@������������������������       �      �<             �?�t�bh�hhK ��h��R�(KKSKK��h �B�  ���-2v?�ߛÖ=�?']P�m��/����?R�+��j�?�9;@��?�����q�?��n����?�d���G=w�v�?�9z=2�?�YC���?3S��˿~|�ʉ����r�:���l�	VB��𿹘el���?H͊�wo�?����g�?84u�w�?�i�'9v?�~�/��?@E0u	��|�C�X�7��]���]H��~66����?�p����%פ�a���ݎ^%ֿp��e�)�?OA�/���j��̦�T�6������;Z�讱?�6�߱K�?��K�3��?�'�1�?�\�鬺���׽����ۅS�T��Yw�֧�����\sAӿrF>Ӿ�\rtu_K�̨�3vu꿺M�R����_�ñ��PG����_�VV�׿�M��z��?�-��K ��_y�5%���̷��ӿ$&S�K�?����M-�?r�� �?J�x��Ŀ8����5��ݨ��鿂�'+Y��?-�F7�	�?!l��HJ�+��C��?�����?� � �@�	u�Q��?�!�ɨ��?%���7�?J�&��?�D��ӳ���u��[���Ao��N�P�ȵ?X*!����?�j��_G�mn7�;���jS:[�⿽��F��D��_��m3 ��0&?�s6�����~��?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KSh�hhK ��h��R�(KKS��h��B(         2                 0�"]?Ko9V�?�           �}@                         ���?*7çg��?\           �u@                        `�[�?�����?;           �s@                        �_D�?�S	!Å?(           �r@                         �Mm�?�pT�ك?'           pr@                        0���?��"��?           �p@������������������������       ��n喜z?�             o@������������������������       �j��IAI�?             6@	       
                 �_W?rr�c���?             9@������������������������       �`,*���?             8@������������������������       �      �<             �?������������������������       �     ��<             �?                        �Q��?؅���*�?             3@                       ����?��V���?             @������������������������       �                     �?                           �?@��@;	l?              @������������������������       �                     �?������������������������       �      �<             �?                        �~��?WL)��,�?             0@                         @��?y���8?             @������������������������       ���b1k?             @������������������������       �      P<             �?                        @@��?t� �z?             &@������������������������       ��ށ\`r?	             "@������������������������       ��">�+�V?              @       #                 �Y�?hP�?!            �@@                         �9��?�'��t?             5@������������������������       �                     �?                         ���?lI&:;�o?             4@                        �R�?�Q�#�f?             ,@������������������������       �                     �?������������������������       ���%���b?             *@!       "                  ���?���,�?o?             @������������������������       � JSl�'?             @������������������������       �@����v?             @$       +                 X�X�?�Rc���?             (@%       (                 @�{�?n��Sy?              @&       '                 `�?��i�p?             @������������������������       ��5���]?             @������������������������       �      P�             �?)       *                 0
��?��n�a^?             @������������������������       ���n�C�#?              @������������������������       �                     �?,       /                 0B��?���V@<?             @-       .                 4�@�? <<(;�>              @������������������������       �                     �?������������������������       �      0<             �?0       1                 �.�? �����>              @������������������������       �                     �?������������������������       �       <             �?3       D                 Э=e?�*�FTk?|             _@4       =                 hJ��?�V��mi?             4@5       :                 ���u?���yj?             &@6       9                  p��?<��'��H?	             "@7       8                 �N�S?���	S?              @������������������������       �                     �?������������������������       � �q
[�>             @������������������������       �      8�             �?;       <                 �ny?͇ �?              @������������������������       �                     �?������������������������       �     �F<             �?>       ?                  ��d�?ȡnN�2 ?	             "@������������������������       �                     �?@       C                  ���?N�	9?              @A       B                  ��? ��wY �>             @������������������������       �                     �?������������������������       � PS��>             @������������������������       �       <             �?E       F                 0r�k?�2@�9�i?h             Z@������������������������       �                     �?G       L                 `�լ?��5<�_h?g            �Y@H       K                 ��ܯ?��h2j?             @I       J                 �\ͥ?���Y3?             @������������������������       � ��� �>              @������������������������       �      0<              @������������������������       �      P�              @M       P                 `�0z?>�O�/�f?a            @X@N       O                  ���?��^ˠ {?             4@������������������������       ��rb7�h?             &@������������������������       ����	�R�?	             "@Q       R                 0���?��}���Y?M            @S@������������������������       �����YjG?             @������������������������       �>\)
pX?H             R@�t�bh�hhK ��h��R�(KKSKK��h �B�  �AKi�C�����U�q��lk#�M꠿a Z��g����-�B��C'�<י�e?��mܿJ��C��?6���p�����~=��e��t)]�i�j���?��$�ձ���*��ֿ8x�K&�鿌j�Y�ܿo��OG��������Q���Џ����w���?���b���?߀�ڇ���q��
��1�t�J������t�F\�?	E6oƵ?V�e:�濕K�^pķ?V�0�s�?�X-�_�?����??\��ޖ�?G�O��?l�8��%�?;B��J���"�4���=�Ae�K��ឦ�Z$ȿ7��\o��^��6!ÿ� 6�E��*�1���F�i����?���<�?�t�Nc�?�w#F�?����Ҧ?�d��k�?�2]�<�?��juߠ?��Y�pC?��T�9_���Ω��"���3��TŚ��Y�5E濇�X����4d,(��?ǚ*�������#�f���Yև�@8Fj��?�i��?
��jIM�?��<+ǡ?F�\���?��� 8"�?4d,(��?bf��*�?���L�? ;�}Q[�?�LC:�ض?b4�ܩ?HQ`=�?Ł��N��?7������?1�1D��?���V��?ے!�s�?h���4ѿ}В �?/�)Q��?��h���?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kch�hhK ��h��R�(KKc��h��B�         2                 �C
T?�mU�>��?�           �}@                        �U���Iwa/~�?U            @U@                         .:q?[��]9�?#            �A@                         e	a?{]p
u�?             ;@                        �$?Z?��̫�ώ?             ,@                         �^��?H�»:{?             &@������������������������       ��h�p�j?
             $@������������������������       �      �<             �?	       
                 �؉�?`���(lA?             @������������������������       �                     �?������������������������       �      P�              @                        ���i?$�\�?             *@                        -�?���p~ݦ?             @������������������������       � mk>e?              @������������������������       �      ��             �?                         ���?�]�%[�?
             $@������������������������       ���2��?             @������������������������       �ԁ��&<R?             @                        U��?���3̐?              @                        �돱?�9���_?             @                        `焘? B���2?             @������������������������       � �vN�4�>              @������������������������       � "s6
f?              @                        ��ǻ?�Z���?              @������������������������       �                     �?������������������������       �      0�             �?                        褍�?ċ�V��?              @������������������������       �                     �?������������������������       �      @�             �?       )                 P^N<?�T�BVx?2             I@       "                 �
OW?�
�U�W_?              @@        !                   ��?�{Ԝ��?              @������������������������       �                     �?������������������������       �                     �?#       &                 0�z?,�|�P?             >@$       %                   ��?8���N?             4@������������������������       �(�KLTJ?             1@������������������������       �������>             @'       (                 Ъ
�?�W�Z�u??
             $@������������������������       �����O�:?             @������������������������       ��bph%?             @*       +                 �:W>?1�=�E�?             2@������������������������       �                     �?,       /                 ����?_�{��H{?             1@-       .                  p<��?b�!��p?             @������������������������       �A}��}f?             @������������������������       �      P�             �?0       1                  ����?W���
y?
             $@������������������������       �����8?             @������������������������       �'C�5��t?             @3       J                 ��_i?�Ⱥ�m�?�           0x@4       ?                 0�W?N��cYJ�?$             B@5       :                 ��l^?�d���o?             ,@6       7                 ���T?H���5J?             @������������������������       �                     �?8       9                  н��?(Rl�F�D?             @������������������������       �  �Y�>              @������������������������       ��p��3�F?             @;       <                  �T?�&�$Gm?             @������������������������       �                     �?=       >                   �x�?��`�T?             @������������������������       � ���+?             @������������������������       �      p<             �?@       G                 �M�h?�xy�̀?             6@A       D                 �F�f?iޗ07}?             4@B       C                 �94W?(h� �~?             .@������������������������       �H��i<}?             @������������������������       ��Zڀ�.t?             &@E       F                 �\8?�p��[a?             @������������������������       �h�]]0�C?              @������������������������       �95�M R?             @H       I                    �?��G�:xn?              @������������������������       �                     �?������������������������       �      @�             �?K       X                 ��_?m��/Q_~?_           �u@L       S                 ��\�?��&1R�~?�            @a@M       P                 �y��?�)����y?�             `@N       O                 �R��?�����?/            �G@������������������������       ��)��}?.             G@������������������������       �      p�             �?Q       R                 ��/�?��ǯT�r?R            �T@������������������������       �Dn2٥,�?             7@������������������������       �{�����b?;            �M@T       U                  @��?�~>�a �?	             "@������������������������       �                     �?V       W                 �!�?a\���S?              @������������������������       �h�w̛J?              @������������������������       �7���:7?             @Y       ^                 �9a�?U�Y�(^}?�            �j@Z       ]                 PY�?3-�o��?             2@[       \                 ��,? �����?             1@������������������������       �                     �?������������������������       �
�|qBy?             0@������������������������       �                     �?_       `                 `~��?�Y��v?�            `h@������������������������       �                     �?a       b                  ��~�?�m��zTu?�            @h@������������������������       �                     �?������������������������       ���S�/t?�             h@�t�bh�hhK ��h��R�(KKcKK��h �B  s*$;��'?9���v��>�J��(���Ǝ�����rc�!@͙�i��r���'!A�������"��������?P�� 7��?�[��C�?�O�`v�Ͽ{�e�����SI��� ?�t��z?я����@;��:�13�HE%�q��碱?��[��@�?-=z� �?���N�?'%w'�?$�>����?h='��I�?B��MZ��?��Z|�|��;���<�`J�	>濗�+C�?H��O��?�W����߂��迌F�\�V�?�-^�+�?)����?��x7+w�?W�k�#�?u���#�?GR�38��?����g��?�������E��K\w�����dYV��Ͱ�k�|������w鿐�)�X�?���k濽%�y_��?̰���r?�� �!�?���C�?v͸yԯ�?]�>�c]�?��y8#��?�S�|��?����E��?a�*��^�?�i0t�?|iZ@���?:K/Ff��?�`R�?`�r6��?@�4��?�n5�ܫ?�(Cd�/Ϳ���ho�?�~�������A� ����vǌ�?�d8�0�?����Ք�?d-���?�5�"h��"4�����pb��a���WA���p�,�ڿ�7R}j�rP]�����"g-�?�� c0ݿ\CK#��?0���!�?gY�sF�?«F����?�%։fο�P�kg�u?�=�Ӳ?�`؍�C�?
b�ex�?�=�����?1�9"�?ɽ^�p+O���4Tk쿬]k}�5?���f,�?z�r2���t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K_h�hhK ��h��R�(KK_��h��B�         (                 ��l?�]a��?�           �}@                        �sM?C(QL�F�?A            @P@                        �j�a?W�~�?             ;@       	                     �?���ƥޅ?             5@                        ��k?�Sp�mj?             @                        ,��??���M�`?             @������������������������       �                     �?������������������������       � ��/���>             @������������������������       �      A<             �?
                        ���U?�j�W�?             0@                        ���L?�D��<�y?
             $@������������������������       �ff���c?             @������������������������       �8���P?             @                         `���?�����a?             @������������������������       �� �ɳ�2?             @������������������������       ��J(�=?             @                        ��V?��m롶?             @                        �2OF?2�[Fn�?             @������������������������       �                     �?                        ���X?.	�\�la?              @������������������������       �                     �?������������������������       �                     �?                        �Ib?@�q����?             @������������������������       �                     �?                        �@�? �q˫a?              @������������������������       �                     �?������������������������       �      �<             �?       %                 а��?@)���ˍ?&             C@       $                  ��M�?�0�h��?$             B@       !                 Ps?�ؙ�a�?#            �A@                         P�kl?M��hm�?             8@������������������������       �tʧ�qJ�?             7@������������������������       �     ��<             �?"       #                 @Ұ�?��u�rv?             &@������������������������       ��@,o?
             $@������������������������       �      d<             �?������������������������       �      ��             �?&       '                 �G�|?�Et@��V?              @������������������������       �                     �?������������������������       �                     �?)       D                 p�v�?,�y"Z*�?�           py@*       9                 �kd1?¨-ۓ�?�            �d@+       2                 �bS?�P��g��?K            �R@,       /                 �U����\��?             >@-       .                  8�1?&�FΪ�?             (@������������������������       ��/m[�?	             "@������������������������       �}>�3I�?             @0       1                 �l?0�E�M?             2@������������������������       �<� z��2?
             $@������������������������       ���$�!�P?              @3       6                 B{�?�%͹�?-            �F@4       5                     �?P�t:o�?"             A@������������������������       �d�V�_�?             @������������������������       �zp���?             =@7       8                 �5W�?�pv�t֏?             &@������������������������       ��#�mt2�?             @������������������������       �l����i?             @:       =                 P��1?H�a�&y?Y            @V@;       <                 Xān?��5[e�B?              @������������������������       �                     �?������������������������       �                     �?>       A                  ��~�?�.�w?W            �U@?       @                 vO��?� �F�z?              @������������������������       �                     �?������������������������       �                     �?B       C                 �~j?��	u?U            @U@������������������������       ��p��V�u?             1@������������������������       �*9��Bs?D             Q@E       T                 �I�?��;ֱ��?�            `n@F       M                 ��6�?N�U��?�            �f@G       J                 @Ws�?���k�?�             f@H       I                 �N��?�]vL��?             &@������������������������       ��qs]�B�?
             $@������������������������       �                     �?K       L                 �7�?a�����?�            �d@������������������������       ���bT��?o            �[@������������������������       ���� �?6             K@N       Q                 �f�?����?             @O       P                 h:��?��U�9�i?             @������������������������       �                     �?������������������������       � �T�x�?              @R       S                 �'�?��p	��!?             @������������������������       �  +X���>              @������������������������       �      �             �?U       Z                 x��?]��B<z?=            �N@V       Y                �톟�?X��]�I�?             @W       X                 �N��?�I���?             @������������������������       ��얅�l?              @������������������������       �                     �?������������������������       �      j<             �?[       \                  ��?b�d!�g?9            �L@������������������������       �                     �?]       ^                  L��?�d!o|�c?8             L@������������������������       ���@�?              @������������������������       �`mt�X?6             K@�t�bh�hhK ��h��R�(KK_KK��h �B�  a�=_��Q?�.���?�ՆQC��?������?�)�J)�?ԏ�$�:�?�;M��L�?�DF]�?��-h���?���љq���z����?��.�|[ݿM=9���?|o�Ն����el1鿨k�O���t����?�����?ss�/��?D�[b�4�?�s�����?��k6^�?��5{a�?�_%��?̺3A�?Ӄ�=� @27I�!@^��ce��C������ub�G����A,���I�y�࿏���G�?����E�?�"��`��?W������)�m<�?� 0�ݺ�?_���L�?jq��ֿ�?�[�=�s���1��5�����{U�}?����D��?wg�.'F�?���ظ��?J/~�������C�K�-���J�a����k��\�\�b������˹��+U'��T��c��?6�%�:�?	2�L�迊�J�X8?�?O���?K�l�L�?�����?��O�d�k�'��e�N¿!)�3���	$ej3���x[� ���?�lڿRx�?���?W}o/�3{?��-�E�?�%�?vַ?���l�R�?�q�ʻJ�?���.�{?@��hљ��k�y��?����S��?Z�qP�?+����c�?_�����?�`1馗���&(�忟��|�5�8��u��t���NRſ���vп���D꿑\�7�_��ۃ�Z�?��Ocp�����^1Dk�?6R���A���Q]���?���bDۿ�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KGh�hhK ��h��R�(KKG��h��B�                          0��?��qg�:u?�           �}@                        �9�?�pf,�J?�             i@                        �i�?S�L��eC?�             i@       	                 �vZ�?E�r̼9?�            `h@                        �6J�?!�)?xk8?�            �g@                        P�~�?x9�u�5?�            �g@������������������������       ��v�2PC1?�             f@������������������������       ���oO:�I?             &@������������������������       �      `�             �?
                          +Y�?`_�����>             @                        쯰�? ����>             @������������������������       � ������>             @������������������������       �      �             �?                        x5W�? `�a�_>              @������������������������       �                     �?������������������������       �      л             �?                           �?j�BaZh?             @                        `ju�?���w�3?              @������������������������       �                     �?������������������������       �                     �?                        �d��?��?ӌ5?             @������������������������       �                     �?                        ��6�?���?���>              @������������������������       �                     �?������������������������       �       <             �?������������������������       �      �<             �?       *                 �k��?dy��fˀ?           �p@       %                 �b'�?RN�}u�?(             D@                        P#��?h�P7[�?%            �B@������������������������       �                     �?       "                  �~��?�=%)B˂?$             B@        !                 �;�?"��XaT`?	             "@������������������������       �@9��U[P?             @������������������������       ��4�r;J&?              @#       $                  �DN?r�O�?             ;@������������������������       ��	�遒?             &@������������������������       ��5���=?             0@&       )                    �?������?             @'       (                p�K=�? hBl�u?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?+       8                   p��?o$Υ��s?�            �l@,       1                 �qҍ?bw���r?�            @i@-       0                 p �?��o�c�v?�            �b@.       /                  �6��?mGg�t?�            �b@������������������������       �q8��[q?�             a@������������������������       �3����?             *@������������������������       �      ��             �?2       5                 �p�?
�$F�CK?4             J@3       4                  9ר?��4KzC?,             F@������������������������       ��v;���[?             (@������������������������       ���'g��?              @@6       7                 �~�?�U1��\?              @������������������������       �                     �?������������������������       ��N�Y�n	?             @9       @                 0�H�?���iis?             =@:       =                 T�Y?���F�d?             &@;       <                 p��?`��!��O?             @������������������������       � �9�FI�>              @������������������������       �                     �?>       ?                 ��L�?�b�a�B?              @������������������������       �                     �?������������������������       ���D�|"?             @A       D                  EC�?%�Xs?             2@B       C                  ����? �*ԓ?              @������������������������       �                     �?������������������������       �                     �?E       F                 �2*�?�d~�D?             0@������������������������       ����0=?             .@������������������������       �      @�             �?�t�b��      h�hhK ��h��R�(KKGKK��h �B8  �i�&:�T�\�k]r���Q�!q및�L^�����%��Œ����WG����)��:�J0ֶ������翕4ق͌?��qmP�?���v��?󹂶��?��m�f(�?�W��b��?�Q�$M��?�]�ݟ1�?hdu3	��?�����?A�h5��?ĭ�^���?�����忀"�W�N�?� �N�?~^T ��?;�}�~��?�z�@�X�?������?p�Ͼ��?��V%��?�︁`�?t��:�7����V	���e%�H�;�?�Y����?'2�}�c�?��D}V�?漢��d�?�= a�r�(�kw�RT�����?Nh"%�@d���gL�wf�p%�{��xP�������H%��/"h5x�����EAP	�b��DgF�"lJ�?F@�>s�?�"٫��?�J�l���?��f���F?'�o'���G�S����?T�����?�M�bi?��z� ��a����j翸xh�!�忚�\�J�?��������C�?�?
Y1�?�$�CNo�??=����?-*�ɑ�?�ȍ����?EiN �m�?��kO���?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KMh�hhK ��h��R�(KKM��h��B�         8                 P�}A?�.Tm�l?�           �}@                        0ϐ? �t?            q@                        83<p?U0M���h?�            �l@       	                  `���?�M83a?W            �U@                         Pmj�?�I<ThT?             @������������������������       �                     �?                        �\�x?��L��C?             @������������������������       ���#�'?             @������������������������       �      @�             �?
                        �x?�\5�_?R            �T@                        �C
T?@?�T?G            �Q@������������������������       ���ؚTI?0             H@������������������������       ��ⱍK�U?             7@                        жd|?���S)bw?             &@������������������������       ���>31g?             @������������������������       �0��$-�d?              @                        ���?N�KtPl?�            �a@                        ��{�?��_�!�l?�             `@                        ��Yk?�n^㰖m?u            @]@������������������������       �,�6�Z	m?U            @U@������������������������       ���Q��j?              @@                        P��?�`7ՇQ?             &@������������������������       �C�S�c�A?             @������������������������       �� �,�8?              @                         �9��?`�$хW?             *@                         �\�?�0h(i�(?             @������������������������       � �7_?�>              @������������������������       � <㣹:?              @                        �:��?M��PI?	             "@������������������������       � ���s�>             @������������������������       �\>�%��?             @        +                 ���?kD��ߋ?,             F@!       &                 �>�?��}"�?             .@"       %                  ���?j���-�{?             (@#       $                 pM�4?ڠ�n׺q?             &@������������������������       �x8c��`?
             $@������������������������       �                     �?������������������������       �                     �?'       (                 @�j�? y�N��?             @������������������������       �                     �?)       *                    �? ��vO�_?              @������������������������       �                     �?������������������������       �      `<             �?,       1                 �� �?#�OW��k?             =@-       .                 P�&�?���m?             ,@������������������������       �                     �?/       0                 �X\�?&�2w��Y?             *@������������������������       �䠪%GR?             (@������������������������       �      P�             �?2       5                 ���?�ގ�E?             .@3       4                   ��?�_>B�@?              @������������������������       �Pu�5A&?             @������������������������       �`ͻ�x1?             @6       7                 ��H�?�����?             @������������������������       �                     �?������������������������       ���ȟ֘?             @9       @                 �0;B?�@�J.fX?�             i@:       ;                  ����?1x��y?             @������������������������       �                     �?<       ?                  ւ�?J �H?             @=       >                 �ig�?��KB�?              @������������������������       �                     �?������������������������       �      �             �?������������������������       �                     �?A       D                 �Q]C?�Bv���T?�            �h@B       C                  ?X�?8���}P?              @������������������������       �                     �?������������������������       �      @<             �?E       F                 ��C?�K��ZzS?�            @h@������������������������       �                     �?G       J                   s��?�l�v`Q?�             h@H       I                   E(�?\/k(��X?=            �N@������������������������       ����c��G?,             F@������������������������       �ﴱ�Gh?             1@K       L                 �j��?r=�YhJ?�            �`@������������������������       ��4�js�i?             3@������������������������       �6�!�1?q            @\@�t�bh�hhK ��h��R�(KKMKK��h �Bh  ��R�lS?&��T���?1Cx�Va?�����y�?^nH����F���!��?Ү����p�S�s濒s��翛/p!��?�gF��?9)��b�?���q��?@�x�I����a��t�b�>��?��T�Au�����怿j���s���_�F˿g-,�?���G��[+�!����p�� S7!\�?T�o����?����6�?��W��?��#R1ux?��g�S�?�MTJ��I�vd��?��ܼɅ�?��<�E�?��:xw�?�/�Z-�?�����j�?4Æ���?�=�s��?b�����?��Ȋ���?� ��?��fS�i�?D2�u2B�}�vw;ɢ?bB�v��迹c4��f�?zKo���?���N�������>�5������ '7��?��%翯��w��;֥�e����"��'z����->�
�&����]�!��1�~񣿃�S�����h4mL{�忪$t�+��|E��r翕8���L{�5�9�?��_)��?&����/�?�}�9�"������OT�{���L�8��]3L�I'ο�^W�5追�E&�vi���5���?  [��޿�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KIh�hhK ��h��R�(KKI��h��B�                          0���?6��Y'�r?�           �}@                         2V�?/+7��Kp?�             m@                         ����?�\d��@o?�             m@                        ���4?\���Hl?�            �k@                        p_Q�?�_�e�Bl?�            �a@                        ���?�%���2o?i            @Z@������������������������       �lxq3�Hi?]            @W@������������������������       �aS:(`pz?             (@	       
                  ��?`��t�[?&             C@������������������������       � F����>              @������������������������       �?��@'Y?$             B@                        �b'�?I�j?P             T@                        �rq?0u�]IZ?<             N@������������������������       ���c�V?"             A@������������������������       �E �B�KY?             :@                        0� K?���P�{?             4@������������������������       �/��S�?
             $@������������������������       ��:�C�FK?
             $@                         @���?H0dP�?	             "@������������������������       �                     �?                        �y���՜��l?              @                        .25Q?8�d�p?             @������������������������       �                     �?������������������������       ���'�P?              @                           �?���?             @������������������������       �p�x��>             @������������������������       �@�����>              @������������������������       �     @�<             �?       0                 0�Z�?BA/��t?�            �m@       )                 P #�?�~�4� j?&             C@       $                  �?h}y��Of?"             A@        #                 P�%�?6+ǉ�(M?             :@!       "                 `��??��
QA?             9@������������������������       �q~7l�@?             *@������������������������       �����e4?             (@������������������������       �      l�             �?%       &                 �Wۘ?�L���Jw?              @������������������������       �                     �?'       (                 `<��?�vnV�g?             @������������������������       ��r��:~L?             @������������������������       ��&3�tS?              @*       +                  �_�?�57��:T?             @������������������������       �                     �?,       /                 �b$�?�o�.�;?             @-       .                 ���Q? O#�1�?              @������������������������       �                     �?������������������������       �      �             �?������������������������       �      �;             �?1       @                 `�C?K��z��u?�             i@2       9                 `�}1?��k?�E�?N            �S@3       6                 �V}?��xŏ�x?D             Q@4       5                    �?�~ν�F`?             @������������������������       � ��mB!?             @������������������������       �      `<             �?7       8                 �ڡ�?Nt�axw?@             P@������������������������       �F���Yq?             8@������������������������       �*�媮x?(             D@:       =                   ���?|^�!��?
             $@;       <                  1��?�Jn��V?             @������������������������       �                     �?������������������������       ���#{M�:?             @>       ?                 ����?؃h�w=�?             @������������������������       �                     �?������������������������       �t��|dw?              @A       B                 ��C?�[ 3�\d?{            �^@������������������������       �                     �?C       F                 �؟a?��V��^`?z            �^@D       E                 0�?p���Jn?!            �@@������������������������       �~��l<�{?             @������������������������       �*:�}*�b?             ;@G       H                    �?��U?�S?Y            @V@������������������������       ���9?)            �D@������������������������       ��_k�[?0             H@�t�bh�hhK ��h��R�(KKIKK��h �BH  ��2�[8��.��OFu?��#�ݪq?�D�e?�]$��\p�l�i�s?�Ё�:������o4I�?����N����:�� �?P���g�.��~�G�?����1r?�v+�IĿ��]���?Y��u�?ܰ��?(����ſ�K�
\�?������?��?	�D}�k�?���I�;�?�[aO%��?
(�����F�Ȣ忌6�k���b����?���VC�w��i0����V/]�z���%i ��훿C*�c헿�R��ˡڿe����L濗���Ba�'�������9���y�0&m���k
���D��A鿈'̝ �?����}�?���U�?���E�?���.�S�?��?���?C�4�hr�;�Pz�B�ΦE�駈��ڔ�dO?�`�i趿Ҡhd��:������%��{?�<��i�?>z
@�¿p��=�����5"���2p�)~�?}-��x濨�'��Rѿ*�����A�RM=�Y��Als{?�fS�M��?"�sI !s?2D�B�?Z�s�NԿ��
��C�?�hT3|f�z_�(k����]�b�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KYh�hhK ��h��R�(KKY��h��Bx         *                 pK�b?n}4��]?�           �}@                        �%�?�:r�Ja?d           @v@                        �)�?��-�0ea?X           �u@       	                 p�O�?o�a,a?R            u@                        P�b�?P�*��]?%           Pr@                        P�$�?0�~��Y?$           @r@������������������������       �]�u~�T?           �p@������������������������       �{PONdr?             5@������������������������       �      ��             �?
                        ��?�~���m?-            �F@                         Pmj�?���TS?             &@������������������������       ��v��>��>             @������������������������       �G��žM?              @                        0��?j���Ho?"             A@������������������������       ��E%~-�N?             <@������������������������       �M����i�?             @                         ���?��2��fb?             @                        �w\�?��t��J?             @                        �)�(?`�K��]?              @������������������������       �                     �?������������������������       �      <             �?                        ^��?x{C6��'?             @������������������������       �                     �?������������������������       � +��Ϸ>              @������������������������       �      @�             �?       #                  ���?�Jp�D?             (@                         ��d�?,���gB?             @                        �'�?Pm�5j	?              @������������������������       �                     �?������������������������       �                     �?       "                 )g�?�m���8?             @        !                  .�?���l\!?             @������������������������       � �+S��>              @������������������������       �       <             �?������������������������       �      $�             �?$       )                �톟�?�@�^(?             @%       (                 tU�L? яDK��>             @&       '                  vb�? M%Ik�>             @������������������������       � ���V�>             @������������������������       �                     �?������������������������       �      ��             �?������������������������       �      �             �?+       >                    �?�ڷ)AH?t             ]@,       /                 ��g?��E�}�4?4             J@-       .                  @?��?t��>��.?              @������������������������       �                     �?������������������������       �      �;             �?0       7                 �C�?Ɖv+�0?2             I@1       4                 ��K�?䮎ȳ�<?             *@2       3                 ��?�L�~�> ?             @������������������������       ��=�p�5?              @������������������������       ��L<���>              @5       6                 @9A�?�=�F�%?	             "@������������������������       � GC6��>             @������������������������       ���x�: ?             @8       ;                 ���?��)�??%            �B@9       :                 �K��?Șv�J?             <@������������������������       ��+3?             :@������������������������       �`3��
�?              @<       =                  z<�? 5��>	             "@������������������������       ��o{u���>              @������������������������       �      �;             �??       N                  �j�?�b� $�P?@             P@@       G                 P���?���|I�U?,             F@A       D                 p��?Р2
�J?&             C@B       C                 0���?H��?�5?             9@������������������������       �2Ū�,?             8@������������������������       �                     �?E       F                 P��?�RF�~NV?             *@������������������������       ������:B?             (@������������������������       �      @<             �?H       K                  ���?��]k:�b?             @I       J                 P�۾? ��7}=?              @������������������������       �                     �?������������������������       �      0<             �?L       M                 �N��?�J���B?             @������������������������       �                     �?������������������������       ���~@�(
?             @O       R                 ��՚? �551�1?             4@P       Q                  �Mm�?�K�6%K?              @������������������������       �                     �?������������������������       �      �             �?S       V                 �B�?<z�y	�?             2@T       U                 �_��?�B����?             @������������������������       ���y� �>              @������������������������       ���* r��>             @W       X                  �g�?��GB�8?             *@������������������������       �                     �?������������������������       �`a�\~�?             (@�t�bh�hhK ��h��R�(KKYKK��h �B�  �\Q�J�H�Nj��r�U�;w�����y�a[��n�D�̓�s��JNoϿ�·0�&�?�
$�'��?AGa�c5��� �?M���/�
���ȶ5�\�3t5��χ�\NeD�9ῴ��G� �?����?�?�H�>6�?0O ��*��h��If�$��@k�(��?�a�h��?&�L��?zV�&=�?M��X
�?{X��M¦?0��id��?�%�G��?�c�D}��?����[��?�>���?M�k�,�?`��.�w�?RR#���?MwV�( �?��z�lQ�?�
�����?Э6j%��?�g-��?�����~�?]�?2�忍��!��?|2_���?RY�C���4w��'濞�j�x����-��?[fڹ�l�?���7�?l���?����?� ��)�?�͢:T��?�a�q6�?�E��a�?�5z�<��?�q[�Z��?�=��<��?�����?=��$���?�-h��g�?�j�(w?
g"R�Q?�4
�1�?|�N��?<$i
�? �XVS��?����F〿�����u?��C�翐�}�Η���[0�
����/�'Q��t� 2翬60p������Qy��3�(�m.�?V�ߊP�?,��+�늿9���TD�"j���?TA�b�?�����K�?+�+=h��?��I�"�?A�
_�?lç��?7�M���?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K?h�hhK ��h��R�(KK?��h��B�         >                  @���?��f�g_S?�           �}@       !                 ��y�?v�f̨S?�           p}@                        ~`��cqA�UL?�            �e@                         W��?��A���]?<             N@                        0S�r?l��.��]?              @@                        0��\?Ҙ��4\W?             :@������������������������       ��ծzkU?             3@������������������������       �Z���˚J?             @	       
                 0)�z?����A?             @������������������������       ��EQ���>             @������������������������       � 0�K�?              @                        ���?�iX��W?             <@                        ��Dm?Xab 7`?             @������������������������       �R�0���S?             @������������������������       � w���?              @                        ��fK?P����E?             6@������������������������       ��V����P?             @������������������������       ��/#�y=?             3@                        ��??�-��[`4?r            �\@                        ЮU?��ag&�1?(             D@                       ���?�٥@
�E?             @������������������������       �                     �?������������������������       �@��fz�>              @                         �~y?0�D��"?%            �B@������������������������       ���x�?             2@������������������������       ��U�ɩ�%?             3@                        ��]?�l�F2?J            �R@                        ��h?���!Q`*?             @������������������������       ��'/15�>              @������������������������       ��ݻC?             @                         H�=R?��0'/?E            @Q@������������������������       ���KSY�M?             @������������������������       ��� ?>             O@"       1                 ��c�?��}%�U?)           �r@#       *                 П�?���1��Y?�            �f@$       '                 ���?4%3�j�^?X             V@%       &                  �A�?���;�o^?M            @S@������������������������       �g��n`V?B            �P@������������������������       ���w�Dn?             &@(       )                   E(�?RhqnrS?             &@������������������������       �                     �?������������������������       �s����;?
             $@+       .                 P^& ?�����R?_            �W@,       -                 �+@?��=)��`?             @������������������������       �                     �?������������������������       ��U�̈dA?             @/       0                 pH'�?m���N?[            �V@������������������������       �D�+#U�J?Z            �V@������������������������       �      ��             �?2       7                  `s�?s�ؤ.K?r            �\@3       6                  `�J�?]����b?             @4       5                 `P�?@�����>              @������������������������       �                     �?������������������������       �      ��             �?������������������������       �                     �?8       ;                 `2�?p@	(��H?o            �[@9       :                 pU�L?���%,i%?             =@������������������������       ��'@r�!?             .@������������������������       ��A�ǥV?             ,@<       =                  �9��?��/N?R            �T@������������������������       �6�>�p�n?              @������������������������       �w.K
iA?J            �R@������������������������       �     ໼             �?�t�bh�hhK ��h��R�(KK?KK��h �B�  �Gq�"�Z��/4b7��4�d��t�U�;%v��Z�?�?|\���>K�����x>������&"h��x�NU9}�?� ��2�?��p��.�?U_�wlc��/��/C��K�濵��4�p�k$���ψ��^�濔a���ڿ���=~�F���9D�\?X�A�����*�2����?,��!N�ֽ)���?��m����?]6����?�hFt�Lu�D��x��*�;�LS��������:��l��Ҫ�;Z߿ �M�ſ����ĸc?m�+�){?�#eR_5�?�Ғ�X
�?J@����?EJw���?�L���:�������|$	�������F��^����D	��|b��l�?���U���^L;�GO?�Ou(�:t���Q���?V`^}�q��j^Ь�?�8=�7�s��
3ƿ��"?�Z�������?��0O�u�:8̨y���y=�a��]v��ޠ�S�~|��[��,]E��?�5y�8�ҿI���?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K=h�hhK ��h��R�(KK=��h��BX                          �$?Z?Ǔ#8x�Y?�           �}@                        ��ϫ?C_��b-[?             ?@                        � �l?J�����S?             =@                        Э�L?4ˎ��N?             8@                        hì+?I����E?             &@                        X��?��X��I?             @������������������������       �h��"*?             @������������������������       ��d�l��F?             @	       
                   �0�?F�%��?             @������������������������       � ���ʆ>              @������������������������       � rtk���>              @                        ��g�?B��"ޒD?             *@                        �o�O?��g��3C?
             $@������������������������       ���� ��+?             @������������������������       ��z�X:�@?             @                         0+Y�?�)��t� ?             @������������������������       �@^�����>              @������������������������       �     ��             �?                        �~�? 
R�{@?             @                        h��a?+�����>              @������������������������       �                     �?������������������������       �      �;             �?                         I��?0ɰ�[K$?             @                        �{�w? �?S��>              @������������������������       �                     �?������������������������       �      �             �?������������������������       �                     �?                        <�vx?��F���Z?              @������������������������       �                     �?������������������������       �                     �?       <                  @���?����zY?�           �{@        -                   �G�?���$"JY?�           �{@!       (                 ���?ҁ��07T?7            �K@"       %                 �%��?�m�T?              @@#       $                 �d�p?�<ǌ�P?             >@������������������������       ���H�3?             @������������������������       ���)���Q?             7@&       '                  ho�?@�8��C?              @������������������������       �                     �?������������������������       �      <             �?)       ,                   ���?��\OO?             7@*       +                 `��?�`D(`�:?             6@������������������������       ��wl��]3?             0@������������������������       �l��|�2?             @������������������������       �                     �?.       5                 �SpR?��Ѳ��Y?�           x@/       2                 ���{?��O��]?:             M@0       1                  �"�?�/��$�P?             ?@������������������������       �;:�nJb`?             @������������������������       ��Q���<E?             <@3       4                 P�,�?0g���c?             ;@������������������������       ��[Nz�g_?             :@������������������������       �      P<             �?6       9                  �P��?Bv8=��X?G           pt@7       8                 �J�?e���� ^?8             L@������������������������       �A)L$�^?             <@������������������������       ��4�a�G?             <@:       ;                 ��_i?��ܓ�FW?           �p@������������������������       �}��L�D?             5@������������������������       ��>�2�W?�            @o@������������������������       �      ~<             �?�t�bh�hhK ��h��R�(KK=KK��h �B�  śO�p:?��QF�?��R]:΄?�"=$��?]-��A�(��dl�*���c#�O:�?M�$I8�࿨��Z��?�*S�߀�?i,�7f��?(����?m�����?Lm����?h�����?q&dT�݈?3,/&^��?�`vh��Q6}ѭ���?���Mv�Q7'�D�忧ZօwX�;�2����{�L�=���Y!q6濉�>���Γ�.���u�-�?ex���?�ƹ��?4Oߡ��E�it,��?����iWq�?dǌ.��V?��.w?U��R�-�?Di���̙��uY	��;���^�S��M.�/��iE�?�j5Lv�?�=��I'�?�X3�����\󼖔�?��a�M_�M�s(+gy?�F�T@|�Uc�,�?vp��$׿��۩c��?+Ir���?j]�@y��T�
|pk����3����ٜTB6�d�U%���?N�ucxU�)gI���⿇\9��d?W.5�x>翔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KGh�hhK ��h��R�(KKG��h��B�         *                 0���?9y �ØC?�           �}@                        P!d�?��3�9�>?R            u@                        @@�?���	�=?C           0t@                        PP��?[?y�W�&?�            �l@                         L��?k���u�$?�            �j@                        ��l�?*g ��/?F            �Q@������������������������       �J�0�/H ?@             P@������������������������       �8ӧ���[?             @	       
                   �g�?AG�k?�             b@������������������������       ��LX��?�            �a@������������������������       �K�n�qSb?             @                        ����?2�7�&�4?             ,@                        �}|�?BX�ظ3?              @������������������������       �T�e|x*?             @������������������������       �      0<             �?                        ��?���7l?             @������������������������       �                     �?������������������������       �U��.c��>             @                        ��[�?�[�Ӽ�Q?^            �W@������������������������       �                     �?                        �aH�>[׫��M?]            @W@������������������������       �                     �?                        �-�?>e��J?\             W@������������������������       �>dda9U?             <@������������������������       ��e��dW@?@             P@       !                 0��?�X�zZ�;?             .@                        �Uq?��a��A?             @������������������������       �                     �?                          �Mm�?ű��?             @                        0>f�?���f���>             @������������������������       �B�l��>             @������������������������       �     ��;             �?������������������������       �      �             �?"       )                 L<<�?`)ٜ_�?              @#       &                 ��'�?pR �m	?             @$       %                     �? ��N@�>             @������������������������       �                     �?������������������������       � @��v>              @'       (                 �ڡ�? K�D^p�>             @������������������������       � �-U@ȷ>             @������������������������       �      <             �?������������������������       �       �             �?+       ,                  ���?46A��L?�            �`@������������������������       �                     �?-       8                 �Q�?�S�>��I?�            �`@.       3                   .p�?��|ÿK?`             X@/       2                  ���?LzS��81?             @0       1                 �b'�?�H?��F!?             @������������������������       ���P���>              @������������������������       �P�ɧ�Z?             @������������������������       �      <             �?4       5                  @?��?��!�K?Z            �V@������������������������       �                     �?6       7                 `���?�f��D?Y            @V@������������������������       �}�Rq�D5?             @������������������������       ��2�Xw�C?T             U@9       @                 ����?4����??%            �B@:       =                 ���?E���j>?             :@;       <                   �0�?�����1?             7@������������������������       ��e�0K)?             .@������������������������       �ͿJ5݋?              @>       ?                 ��Q�?�<jػ�@?             @������������������������       ��8�;K�?              @������������������������       �      &<             �?A       D                 ���?d�	���$?             &@B       C                 X)ɢ?���s��>              @������������������������       �                     �?������������������������       �                     �?E       F                 `���?oV� ���>	             "@������������������������       �:��\���>              @������������������������       �      �;             �?�t�bh�hhK ��h��R�(KKGKK��h �B8  �ի_�0��:�ܶd�1���9�Y��#@i�
o�ã�'�r�����sWW�/ɠQB��C��N��?���D
�w�ks�2h�㿚Ti+��{��=��w?���f��?�Q$�*��?�.��TT�?1����W{��T��w��.�
���ۿ�r��,o?WFL³�?!���-Sc?��>���?_��K��T?�����?p��Uƿ1��򟵕�S(pǂ�H����濫��=?2����d0q�J ��y� �4!B_�?r��_���?�]�W�>��N�!�(���������{���':�j,~f(��n�-�S���zqj�忨%������Ei�f��s4��u?mς��H�?$���cr?-+C�^�?�-����f18~W酿
r!�����$��Y�Ϳ��D��O��G\�4��?�@.>A�?z�T�V��?B	4a@�irf���?����/y��}���q����[JG���p�U�3���*�)s�?[�w��è�]0�������ַ���co�?�� �U��?���k��?���/�*�?�ݮ9dr?L�A}̮�?H��`���?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KSh�hhK ��h��R�(KKS��h��B(         0                    �?�e��58A?�           �}@                        �7d�?��l�UjB?�            @o@                        �n��?�1BD?�            @k@                        �v��?�F�؃�A?�             i@                         �~��?�	,�?A?�            �h@                          s��?ի�^SC?T             U@������������������������       ��B���>?R            �T@������������������������       �p� �^?              @	       
                   ��?����>?q            @\@������������������������       �����K?             1@������������������������       ��Q�b�7?`             X@                       ��G��?5� ��C?             @������������������������       �                     �?                        ��K�?X	�ߜ>)?              @������������������������       �                     �?������������������������       �      �             �?                        0+�?��۷��V?             2@������������������������       �                     �?                         PV��?6
��nM4?             1@                        `��?�����\E?             @������������������������       ���Q(m�>              @������������������������       �                     �?                         @���?�˘�Vg?             ,@������������������������       �:"x3`��>             *@������������������������       �      �             �?       '                 ���@?v�<��?              @@                         ���?$r���Y/?              @                        ��M�?�j��D$?             @������������������������       �                     �?                        ��K�?P�P�q?             @������������������������       � �s �`�>              @������������������������       �       �             �?!       $                  �E�?иB����>             @"       #                �톟�?�6� �>              @������������������������       �                     �?������������������������       �      �;             �?%       &                 ����?�_0?w��>              @������������������������       �                     �?������������������������       �      �;             �?(       +                 ��?r�1��>             8@)       *                 p2+�?��}τ?              @������������������������       �                     �?������������������������       �      Ȼ             �?,       /                   ��?}[0Q�>             6@-       .                  �3��?�c5m��>             5@������������������������       ��?)j��>              @������������������������       �b���>��>             3@������������������������       �      �;             �?1       6                 0�!�? 8Pt�*??�            �k@2       3                  Џ~�?��*���W?             @������������������������       �                     �?4       5                �^B�.?�����)5?              @������������������������       �                     �?������������������������       �                     �?7       F                 p�~�?���aS=?�            `k@8       ?                 ��ҥ?�nw��sC?[            �V@9       <                 ��?�*/&�A?D             Q@:       ;                  `���?H��uЬA?"             A@������������������������       ��p<��F?              @������������������������       ��}ռ:=?              @@=       >                 0)��?[iBcS�??"             A@������������������������       ��4fd=�Q?             @������������������������       �+8�0A,?             =@@       C                  �9��?N�'�aOE?             7@A       B                 �R�־�_��h"?              @������������������������       ���<�O?              @������������������������       ��>����?             @D       E                 p=�?�~�F?             .@������������������������       ����S�E?             &@������������������������       ��o���>             @G       L                 @({�?�l�A�5?�             `@H       K                 г��?.�ޟ��4?8             L@I       J                 @��?���++?7            �K@������������������������       ��D���1?             @������������������������       ���n�&?3            �I@������������������������       �                     �?M       P                 �Y8�?Jk2���3?H             R@N       O                  bB?�֮L�a8?             :@������������������������       ��e���7?             &@������������������������       ��B�	>�>             .@Q       R                  �%�?��:5�'?.             G@������������������������       ��:P�@?             @������������������������       �PB��?*             E@�t�bh�hhK ��h��R�(KKSKK��h �B�  ��x�k@�J/��<W?�a��od?c��E��X?��V[�QR?��f}�g���u�گ�R�[�����b�p?�@]U�A�?�=}ly �?�s����?^�MIi�h�߸��?�g�s��?g�VЗ��?��,�?4݊���?RfT1v?@<���?���&���?x1Y)���?fU�&k9?ϸ<��p忽��&�?�w�;h7x�{z�n|���nğJ��?%P�u���T�ǃ����"��G��Q���zWddAw��.��W��r��	�y忮�;œ�^-e~2�c���i忇��=�[�D���4^����eU���L�Ζ��z:Aa�o�5q��S�X����O�>��Rg��塄\����\�x��(����e��P������+{�P翥t /�΄�;}�4S��?�(˽g��x�i$�+b�`W"=P?�����oa��L��N�}�o�6�K��ru��˿�]#��Ph?��i�UG�?b\Z�:��(}�"ۄ?�g����}�Do&�����l��j̿j��V���?�R)���?-1ݙ���ܳ�hr���Tl����L���oCba�'�UL˨^�%�o��k�U��^�^A����{[��?��p}�9�?C{5��M;�4��x��j��s]��Q�Y�ܿ�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kih�hhK ��h��R�(KKi��h��B�         >                  �~��?�x/x�I?�           �}@       !                  �P��?T��7�E?�            �g@                          �G�? ]�^>?�            �a@                        0.��?my���??@             P@                        �q
�?��OgA?6             K@                        P]ڒ?��(�B?,             F@������������������������       ����RZ=?%            �B@������������������������       � 1%FWL?             @	       
                 �{N? ��Ґ/?
             $@������������������������       ���ќa_ ?             @������������������������       ��c�mhj?             @                        ��?�$,�2?
             $@                        ��w�?!	��	?             @������������������������       �                     �?������������������������       ��p��il�>             @                        pRh�?4|�hZ?             @������������������������       � �_	�/�>             @������������������������       �:`J����>              @                         bB?����`�;?L             S@                        0��\?��e�;?7            �K@                        �U���p3����9?"             A@������������������������       �Mw찉TA?             1@������������������������       ���(sM"?             1@                        �&\?�.�a,7?             5@������������������������       �`V��m?             @������������������������       �">7��54?             2@                        ���p?�g��.�0?             5@                         vpe?m\���&?             *@������������������������       �h���U?             (@������������������������       �                     �?                         0�:�?��*?              @������������������������       �                     �?������������������������       �\;���%?             @"       1                 �-�?����hgQ?0             H@#       *                 n��W?�R�w��U?             ?@$       '                 )�`f?�#�2��Y?             .@%       &                   \��?�¼Ͷ-T?              @������������������������       �ֹ��IR?             @������������������������       ��{-?             @(       )                  �g<�?�|�.tQ?             @������������������������       �<���C?             @������������������������       ���;UD?             @+       .                 ��Ҧ?�
���=H?             0@,       -                 Z��?A0Y�86A?             &@������������������������       ��hS^�2?              @������������������������       � 
=
p�>             @/       0                 ����?ߢ/�pJ?             @������������������������       ���7"u�?              @������������������������       �������>             @2       7                 0I��?Hq̞�6?             1@3       6                   s��?��^!�!?              @4       5                   \��?7!��d�?             @������������������������       � �:�S�>              @������������������������       �9R$�?             @������������������������       �      �             �?8       ;                 ��x�?+�p�З7?	             "@9       :                  4�? ��nW ?             @������������������������       �                     �?������������������������       � �����>              @<       =                �Y�x�?܉�3�e3?             @������������������������       �L!�U?             @������������������������       �|M���&?             @?       R                 `�[�?�gLsSK?           �q@@       O                 `��?��8׋pJ?�            �j@A       H                 �/�?�Bړ��G?�            @j@B       E                 P��?=h�b��F?�             i@C       D                 ��?�u��7:F?�            �h@������������������������       �~G�~�B?J            �R@������������������������       �u�\�ʬG?}            @_@F       G                  ��?$L��#�4?              @������������������������       �                     �?������������������������       �                     �?I       L                 ��2�?OJf��^P?	             "@J       K                 �5W�?��'
45?             @������������������������       ��6��I-?             @������������������������       �      �             �?M       N                 ��O�? ��cJ?             @������������������������       �                     �?������������������������       ���ټ/?             @P       Q                ��Sl�?��Wk�]?              @������������������������       �                     �?������������������������       �                     �?S       \                 �%��?KX-y�_L?H             R@T       [                 0㒲? +$�ro?             @U       X                 �n�S?e�{�WF?             @V       W                  `���? �>�zt�>              @������������������������       �                     �?������������������������       �      �             �?Y       Z                ����?`�f2vX�>             @������������������������       �`�EH�Υ>              @������������������������       �      л             �?������������������������       �      P�             �?]       d                  (��?�.䎺>?B            �P@^       a                 �	I�?�8�2{�I?!            �@@_       `                 p'v�?��_��A?             :@������������������������       ��j��
?             4@������������������������       �$A��
�R?             @b       c                 0".�?�'@�G?             @������������������������       ��C� [�?             @������������������������       �P�\���8?             @e       f                 0���?j4wd�?!            �@@������������������������       �                     �?g       h                 ���?�y�[*� ?              @@������������������������       ���		�?             ,@������������������������       ���e����>             2@�t�bh�hhK ��h��R�(KKiKK��h �BH  ��HQ��C?��8�|n?G�9�M�E?0U|?��s?FP�t|?�0�9�Yr?���1���?�c=���ۿ��O`?��?�G�F{�?�2@����?z&.P�x��#��rt?N�u���n��p$�?�4[5ب��1��º�lVD_~n忦�{�Qg�^{�D$�|�Ӭ1M@ˈ���?��࿪���><ѿ4D��{KU?\����?�����������a�?6��"N�?8�Y�Τ�?���d��?���HWf�A��~���1Uċ�?%���?�kj����?��%���?$�Ѹ{̍?��Z���?�k&Qҿǵ��j)�?��~�:��?�����`�?hz?���I�MS�P"�e���=�����?:zߟ��?���H��?7}�Qx��?�ew� L?�/�Bt��P��p���n�����"��տf���V�忪���ZS�?K��S���?��,���?�����?E����EG?�L#3����,ϛ��?>�g���W��l*cNsl���"|3ie�$�/?e\�-���;a��7a��?����?�ſ�� ��?/�-���?P������?;f!�-Ж��Q�i����S��g�:�z��?�1Ӏn���T�V�f�]d�'���-+�������]��{�|�����W?cor?P%i�?�|��䓏? �V�#�?��J5|�?l�{�K�?�P[z|w���@��k��	�����nޝ���?��]ۤS?�$H]s�?�L�vRR?���k��ګ8��?:��cp�?Npn�?͠�ܼ�?�p��y�!_�c,��?�W/�Z�{�����忍��2�v忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kah�hhK ��h��R�(KKa��h��B8         >                 �6Sz?L��@�3?�           �}@       !                   p��?���3� 5?           �w@                        �,$i?yt�p�3?[           �u@                        �U���|�	�r*?�            @j@                        P�)�?��Ŋ =5?b            �X@                        @aݨ?r_%h�_�>8             L@������������������������       ��#�����>7            �K@������������������������       �      <             �?	       
                   .p�?,����D?*             E@������������������������       �O7�3Q'?             (@������������������������       ����X2�E?             >@                         NA�?d0��_�?p             \@                        ��+a?����cT?i            @Z@������������������������       �\Ξ���>e            @Y@������������������������       ���iҘ�1?             @                         �6��?l��~��,?             @������������������������       �����v?             @������������������������       � BV��=�>              @                         �6��?�i�a9=?�             a@                        �D��>�P�r�6?~            �_@                        ����?���p??            �O@������������������������       �:��E@�>             >@������������������������       ��{�yI�!?!            �@@                        pb�?Zt#\�B??            �O@������������������������       �z��X.?'            �C@������������������������       �9��.�P?             8@                        @��?�����T?             &@                          B�?�B
��	'?	             "@������������������������       �                     �?������������������������       �@(���-?              @                         ��T�?��!��`?              @������������������������       �                     �?������������������������       �       �             �?"       1                 �r>�?����=;?$             B@#       *                 P�bf?1y�
�9?             3@$       '                 �t�?6 ���3?             &@%       &                 ,OF�?�L���>�>             @������������������������       ���J�q*j>             @������������������������       �      �;             �?(       )                 :��?�Y���1?             @������������������������       �                     �?������������������������       �8׽�y
?             @+       .                 ���?��h� &?              @,       -                 �_��?�x�u=B�>             @������������������������       �hO��:�>              @������������������������       �H7����>              @/       0                 ��ǻ?��6��?             @������������������������       �                     �?������������������������       �����?             @2       7                 �%�?[���6�1?             1@3       6                 �o��?��+;$dA?             @4       5                  ����? �S��;�>              @������������������������       �                     �?������������������������       �       �             �?������������������������       �     `3<             �?8       ;                 0A�?p�&r�?             ,@9       :                 �\͵?�>��)�>             @������������������������       �                     �?������������������������       � x��F~�>              @<       =                 ��C�? �A�k
�>             &@������������������������       � ���8�>              @������������������������       �`M)P���>	             "@?       V                  ��?�⭡�k ?Y            @V@@       I                 ����?�
KU?7            �K@A       B                 ��? 0H�h?              @������������������������       �                     �?C       F                  ��^�?$ì���>             @D       E                 ���? �����>             @������������������������       � �e�fY�>             @������������������������       �      �;             �?G       H                  �h�? �oѽ��>             @������������������������       �  �pQ�>              @������������������������       �      л             �?J       Q                 �5=�?�q�@�	?/            �G@K       N                 `���?�����D?,             F@L       M                 @9A�?��%;� ?%            �B@������������������������       ���ȁy�>             8@������������������������       ��4��JY?             *@O       P                  ��^�?�w f]\?             @������������������������       ��CF���>             @������������������������       � �(J]��>              @R       U                  �6��?�{���_�>             @S       T                 �.7�? �dtn�>              @������������������������       �                     �?������������������������       �      �             �?������������������������       �      �             �?W       X                 � �?b�����*?"             A@������������������������       �                     �?Y       Z                 ���?�ɠ1�>!            �@@������������������������       �                     �?[       ^                 �٠�?���R��>              @@\       ]                 0���?�����?             @������������������������       � ���sr>             @������������������������       �                     �?_       `                  �Ȕ?���e��>             <@������������������������       �                     �?������������������������       �l�f�B�>             ;@�t�bh�hhK ��h��R�(KKaKK��h �B  ��P�J�G�$�S��B�
�`�%
>P����v��6n?���c�� �ϡt�UV+�Ʃ�?����C��?���2�ѿq=��*��?���qj��Ɔ��`����n��c\�{��?
i��Qʖ��)y�Ӱ�%�pR�f��su���f_\�o���8��.5�%�'�$=��Q俧�#Ұ��>�/X��Կp��%��?��	ԉF���
��a��E�<濅��1?Aٿ/ӹ(�J��w��\�������2�m5Q}?l����TV�)~�$
ȇ�R���,K�!�闪X���0d��Z�6������.�� ���U���^��?�b��[e?y��J��?����c�`:�af�?��\�-�?G��,��?��R��?+0̗A��?г��լ?YƵTՍ�?�C1�Ũ�?�c<%�?�F�l�?��HC�a�?ٿ�(q��?�JS��?�\cS�~?J�Dr���?�X�a{�?Ŀ���r?*�lכ}?��؊�)�?`j�i�? 4+�x��?�[��-�?Ϊ�]��?�����?kS��Y�?�JT�¡�?0u&���?�y�Eax?�@��v?}�s1��r?�÷L���?_���x�?�Ohxm;�?t5���?�y���?����F�? y��?݊C��?���@m��?�B�/R��?�>nz6?�L�������f?���l&��?ڳ�°�b?.�]%tf�`�'�Je�?o,��忒�҂�h?�6�F���?!H3m*g�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kgh�hhK ��h��R�(KKg��h��B�         2                 0'Fx?Fӏ��,?�           �}@                        ��{s?s�Ͼ�/?h             Z@                        O�z?Ɠ8�/?U            @U@                        �><r?o;r��N+?O            �S@                        @�K?GL{�5�,?9            �L@                        P.�?�� �U�&?             =@������������������������       ��&��j"?             6@������������������������       ����;/�!?             @	       
                 P%�o?^�g.M])?             <@������������������������       � ND.o#?             ;@������������������������       �                     �?                        �0Le?=�����"?             6@                        ���`?թ���"?             &@������������������������       ���ro?	             "@������������������������       � -�TA�>              @                        0p�:?�C��)?             &@������������������������       ���֯?             @������������������������       �
���F�>             @                            �?0�ɦ�e>?             @                        0ꀄ?�'�a��?              @������������������������       �                     �?������������������������       �       <             �?                             ���� p?             @                        ب��? 0�z4�f>              @������������������������       �                     �?������������������������       �      л             �?                          .p�?�:;2�I?              @������������������������       �                     �?������������������������       �                     �?       )                 ،&a?�:�&?             3@       $                 h��@?ܹ֛H?	             "@        #                 ��
w?(mY��U�>             @!       "                  �P��?��19�L�>              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �;             �?%       (                 ��h7?`hz��?             @&       '                 �`>`? �Ex���>             @������������������������       � �4��>             @������������������������       �����i��>              @������������������������       �      ��             �?*       -                   ���?��w0<�?
             $@+       ,                 @��?4��sH��>              @������������������������       �                     �?������������������������       �      �;             �?.       /                  ���?�pkX$
?              @������������������������       �                     �?0       1                 �2OF?�5�%υ�>             @������������������������       �6)�$���>             @������������������������       �`޾��~�>              @3       J                 `ӄ�>���U�Z+?p            w@4       ?                    �?Z!sL_�4?             1@5       :                 ��!�>μC(t`6?             &@6       9                �3�.s?sN�tYy#?             @7       8                 �_[�?)�%=��	?             @������������������������       ���[Į
�>             @������������������������       �      �;             �?������������������������       �                     �?;       <                 P�?*�k퐗6?             @������������������������       �                     �?=       >                 I�@?�Q��~?             @������������������������       �� �G~�>             @������������������������       �       �             �?@       C                   �P�?�q��?             @A       B                  ���>�ezWA�>              @������������������������       �                     �?������������������������       �                     �?D       G                  �Ԧ�?,J��Q?             @E       F                 �m۶? $7;���>              @������������������������       �                     �?������������������������       �      �             �?H       I                 W�h�?���%��>              @������������������������       �                     �?������������������������       �                     �?K       X                 �HM?ϝ�s)Y*?_           �u@L       S                 Lg? m��>L5?             1@M       P                    �?���.Z��>             @N       O                 �vg?�NJ$��>             @������������������������       �t���H��>              @������������������������       �                     �?Q       R                  @?��?}a�a}u�>             @������������������������       ��P�\ �>              @������������������������       ������>              @T       W                 ���I?���25?
             $@U       V                 �  )?��Z�+?	             "@������������������������       �p�ɕ>/?              @������������������������       ��_8��>             @������������������������       �      8<             �?Y       `                 Ш��?�*��x�(?N           �t@Z       ]                 Xbp?L�Z )?�             e@[       \                 p��?�)��2?V            �U@������������������������       �u���z�=?.             G@������������������������       ��ɠIB?(             D@^       _                 z�?�P��/?S            �T@������������������������       �2�,��?             &@������������������������       �k�	��?H             R@a       d                 ��?��a]
(?�            �d@b       c                 ��{�?z6�7"j2?8             L@������������������������       �\?j��l6?!            �@@������������������������       �v��?             7@e       f                 ��Ĳ?����UY?m            @[@������������������������       �*�6��?6             K@������������������������       ���2ҝ?7            �K@�t�bh�hhK ��h��R�(KKgKK��h �B8  �tnú�!�$%- o-g?&2�߳Q?�����?̐D���`?3X�@m�n���A������G��⿭������?+s����?�X�G�V�?�����u�C��?M?ûZI Rӿ��ڟ��?���膿Z�X	��忏�Z����1{ti@+�?���Sx�?�vV ��?pP$�t�?��W�ҁR?�JI*څ?q����?+&	�a��?�TI��9����w�c��z�����d�z *х?��<��?+u�/~?��ifz�?z�b��?A�$��?s�c ?i�?K�3��O�?���U �?�V�D��?(��!(��?��К�?�� ��fe?�<�WK���������i��~s�gc�҅x?���t"��?�,�:q?FFP�a�?��o��b�y<�O����A�x?lSGb�?Ǘ�/ae?�<+9E�`��6?�?R	Ϟ忚Ivc���?�o@#���?�)R�á�?2=��?��/��?�V�¦��?i��h�@u��^�s?6��0�V�X��S��??�i�ׄ��LQ�A���t'([S��jq������b�kwp�/:���{�&��x�Z�s8�3~[U�<jV�q����f�Oe?U�.7��x?�C���i�?2٤!w��?�g;-a?u%���f�?6�p�wh�:sҽˑ�����x���9_�K:T濧��7��"���o���-�v��J�U��3KXd�F����q��@�G��׿���oe�? G
�B�ď���G�?�|��e�ӿ��*,�L?V����w?D	 W֬?	���}4�?4pGR�Y�b��j�ڿ���uQ�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KWh�hhK ��h��R�(KKW��h��B         2                 ��'|?��q�3?�           �}@                        ��{s?�~�Cgx0?w            �]@                        O�z?y�oө1?U            @U@                        �><r?�:1�I�/?O            �S@                        @�K?���mj/?9            �L@                        P.�?�V6Tj(?             =@������������������������       �|�~-#?             6@������������������������       ���
Y�E$?             @	       
                 P%�o?���ȈR-?             <@������������������������       ��)�~�'?             ;@������������������������       �      B<             �?                        �Jh?�>�)?             6@                        ���`?���w�� ?             (@������������������������       �l�1#�L?	             "@������������������������       �zs3�9�"?             @                        Њ�(?&�X��$?
             $@������������������������       ��჆�`#?             @������������������������       ���k�M?             @                            �?���6f;?             @                        P�J?`�笶
?              @������������������������       �                     �?������������������������       �                     �?                        �t�?��Ͻ�?             @                         �JV�?^���SY�>             @������������������������       �                     �?������������������������       � �2����>              @������������������������       �                     �?       '                 `�F�?غ�T�%?"             A@       "                 �R�*?C�� ?             9@       !                  `<��?�s����?             .@                         ��h7?�ͫ��?             ,@������������������������       ��{���?             @������������������������       ��z5�/�>              @������������������������       �       <             �?#       $                  �Ԧ�?(oB��?
             $@������������������������       �                     �?%       &                 �݂�>�5�؀_?	             "@������������������������       �@]?���>              @������������������������       ��3m�2e�>             @(       -                 @u�x?�u�Ѹ�?	             "@)       *                  p�{�?b���2�?             @������������������������       �                     �?+       ,                 ��G�?�i�����>             @������������������������       � &��EN�>             @������������������������       ��dUI�B�>              @.       1                    �?��~�X�>             @/       0                 @ۆy?  ��i>              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �;             �?3       :                 0h�~?8�8�n�3?a           v@4       9                 ����?C%X�8?             @5       6                 �n|?@����#?             @������������������������       �                     �?7       8                    �? �{EI?              @������������������������       �                     �?������������������������       �      �             �?������������������������       �       �             �?;       J                 ���?�b�&3?]           �u@<       C                 �Y�b?�B�@�6?             8@=       @                  V�>&.�[43?             *@>       ?                 �.��? dv`��#?             @������������������������       ��_�@,��>             @������������������������       �       <             �?A       B                 ����?�*�i� *?	             "@������������������������       ��хr/ ?             @������������������������       ���vt�?             @D       G                 ��{�?ر�懜,?             &@E       F                 *\?l�:O�>              @������������������������       ��U�1o�>             @������������������������       ��c��I�>             @H       I                 �Wci?<P����?             @������������������������       �`�)y���>              @������������������������       �      <             �?K       R                 P.�?ܳ�%f�2?E           Pt@L       O                 �\͵?���B�*?             0@M       N                 (l�V?�����>	             "@������������������������       ����R��>              @������������������������       �      �;             �?P       Q                 �u�>�=a�@0?             @������������������������       �                     �?������������������������       �0��w�>             @S       T                 Ѕ !?����2?5           Ps@������������������������       �                     �?U       V                 �<�?�G��ͭ1?4           @s@������������������������       ��̋��b??G            �Q@������������������������       �F����*?�            �m@�t�bh�hhK ��h��R�(KKWKK��h �B�  Ujb�7?����a����� ?�g� S?j�����T�zq}?~�r?.��c@�?���+�
�?	R��}�kP���տp.G)�P濖u�K�~?�Ф�C?آ�&��?o�
�r޿��r�F�?�Hdwu�?}~�E���?��Y 닿f!P��"��-�R�
��9�v_�"��W�I�[NX
h�y����wW��x��+��c��*{��?�kN�s������r���pb�
^����S}�$��0Qv'l�������c���Щ�#�w��u����eHn~�k��C�)����_[����g�˱~Kg?��2�\2a����Y���?�R1���x�_M�K�l�Z�g�����Y�k��?�}C���?�A�$x��? ���?����&z�?��~cݡS?��r�G��?������?���o�i�?0��4��?�c��?��z����?��C�:��?aܲ#>�L?K�,���}?^�3�5�?��U�&�?��3���?#����{�?y;6r��?�͂W�f˿� (1��?m��wg�M�I�U���@�����'}Ww�0�ܵ�?=��;��?�F�O=�?�r�y}�:?����m���މ�&C�u��;��῞��-��?��?gT&����އ��q�&�o���O�Q8�L?�`����?6�A��E?A�Xk��?I��p]���t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KKh�hhK ��h��R�(KKK��h��Bh         4                 �)�?'Ȫ_(?�           �}@                        �6Sz?9���:?�           �|@                        �f��?��nl�$?v           `w@                        ����?[��|N?e           Pv@                        ��?|���?�            �k@                        ���?﵎E�B?�            `c@������������������������       �q,�.s?�            @a@������������������������       �����.?             1@	       
                 ���N?���:�$?A            @P@������������������������       �˸F�( ?#            �A@������������������������       �H����'?             >@                        P�$�?�r�G��?�             a@                        @�P�?lYf��)?f            �Y@������������������������       �
�3ks?_            �W@������������������������       ���K��>             @                        �/��?(�0)'?#            �A@������������������������       �N�E���@?             @������������������������       ��'I�d?             =@                        ���?��J�`�*?             1@������������������������       �                     �?                        ����?�݆��R!?             0@                        PUٰ?��a��?             &@������������������������       �num�Б�>             @������������������������       � HP?�?             @                         ]�?fkU��	?             @������������������������       �                     �?������������������������       �;�e��>             @       )                 �ħ?U@H�Jz�>U            @U@       "                 �C�?T� # ��>$             B@                        XFe�?�
�2-1�>             @������������������������       �                     �?        !                 PQ�? o�j��>             @������������������������       � |�v�c>              @������������������������       � (��lV>              @#       &                 ����?@ВX��>             ?@$       %                 �r��?�<8�գ�>             0@������������������������       ���ʜ�w�>             ,@������������������������       ��U8ln��>              @'       (                 @Ws�?� ��5��>             .@������������������������       �| bh���>              @������������������������       ���c!��>             @*       -                 �H�?�Sg�?1            �H@+       ,                 �\��?@�s4��4?              @������������������������       �                     �?������������������������       �                     �?.       1                  Ja�?�WV1��>/            �G@/       0                 @t�?�r�Ld�>             @������������������������       �@���>             @������������������������       ���"�r>             @2       3                 �2T�?�����>)            �D@������������������������       �                     �?������������������������       �28jv��>(             D@5       6                 �Q�?�;=�6�$?             *@������������������������       �                     �?7       @                 ����?��a�?`?             (@8       ;                  @V��?H�~���>             @9       :                 H�}�? ��UP�>              @������������������������       �                     �?������������������������       �      �;             �?<       =                 ��?`�C�ܽ�>             @������������������������       �                     �?>       ?                 8n��?��AТ�>              @������������������������       �                     �?������������������������       �                     �?A       D                 �D��B��wB�>             @B       C                 �h��?�t�S���>              @������������������������       �                     �?������������������������       �      ��             �?E       H                 ���?�$K�p��>             @F       G                  �1�?�N�|�6�>             @������������������������       �                     �?������������������������       �c����>              @I       J                 �fa�?��&hd�t>              @������������������������       �                     �?������������������������       �                     �?�t�b�1     h�hhK ��h��R�(KKKKK��h �BX  �6f�,���I�q�;�Ф�0N�go's�~D����[�
'?�OW-�T�K����Ŀ1$uV!�׿@�'b�m?�����?��?��i�T_�o�˥j�]3=�A"�?v�?H'�hXX`?��8���?��2C_���@�7}�3e��G�2����'t���PɃj��n��8/ۿ0`���忴Fߐ��t?@��9ٻ�?�s���?�0�f�\?�}#Vm?�W#��{{?6�Kft^�?�߽ǿR�?q)F n��?�2X@z�?[����3i?��5�%`?�t�Z|_�?����iz�?��'vq?!W��i�?]*Z�|�?kF[h�';?<���b���^��Z�?+=2�f�ۂ��R?=	\�ss?_;�g~�?,�.a�?x��B�D?`��Aۋ���P���?[5ީ}?���JT�?�R!�?Op?��X��p�?�~*	ӂ�?$���?�ݗ��?��`"x?䚈6uf�?�U;��}?d e����?_{8�v�?�W�V��3��v��]s��K�/����SH|]����X?S�
!�2A?�:�KS]�?���g��? ���g?	��ߔc�?�A�F�f�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KUh�hhK ��h��R�(KKU��h��B�         (                 )DW?��Q:�l?�           �}@                        p��C?b��	3=?b            �X@                        P���>T�9lM?]            @W@       	                 ��>m?������?             ,@                        �$I�?Z�[���?             @������������������������       �                     �?                         �vg?h��W�>             @������������������������       � ��(Nf�>             @������������������������       �       �             �?
                        ��a?�I��K��>             @                         `���?0�����>             @������������������������       � 9�� �>              @������������������������       �      �;             �?                           �?��Nm��>             @������������������������       �e\��o��>              @������������������������       � �E�@A7>              @                        ���L?�`�I?O            �S@                         DM<?�L���r0?             @                           �?mg<|��>             @������������������������       �H0���%�>              @������������������������       �      л             �?                        x5W�?`v��%�>              @������������������������       �                     �?������������������������       �                     �?                        �x?/�B�܇?J            �R@                        �s�Q?�%�h��??            �O@������������������������       ��Ş>��>             @������������������������       �ոi��?;            �M@                        ��Ɲ?��D��?             &@������������������������       �z���\L?	             "@������������������������       � wC���>              @        #                  p���?�yA�?             @!       "                 �)�H? ��Dih>              @������������������������       �                     �?������������������������       �       �             �?$       %                 (�!�? ��8�C�>             @������������������������       �                     �?&       '                  ����?Ѐfy�s�>              @������������������������       �                     �?������������������������       �                     �?)       B                 вeh?��=�$�?v           `w@*       3                 :F?t<�'B�"?�            �b@+       ,                 �?�N��l?             0@������������������������       �                     �?-       0                 ��lw?4d�K�s?             .@.       /                 @��?p�G�}�>             @������������������������       �`��n�>             @������������������������       ���Q�N�>              @1       2                 �Z�?�t+�j?	             "@������������������������       �fS��P�>             @������������������������       �Z�Q��?             @4       ;                  �P��?5�WFv"?�            �`@5       8                 `�h'?&��`��)?)            �D@6       7                 �r�?�R��]5?             5@������������������������       �&��
o8?             *@������������������������       �#%+�YS?              @9       :                  �9��?��n��5�>             4@������������������������       ��O���s�>             2@������������������������       �,Xy�g�>              @<       ?                 �F�f?�ϟ�'?\             W@=       >                 @+{�?�p�K��?             @������������������������       ���.��U�>              @������������������������       ��F��H?             @@       A                 P�Y�?����2?V            �U@������������������������       ���(?@3?             @������������������������       ����~�l?P             T@C       L                 P\?����r?�             l@D       K                 `S[?��~i�$?v            �]@E       H                 `��?�f A�� ?u            @]@F       G                 `s5�?�A3NsY?             @������������������������       ��?���>              @������������������������       ��	֌R�>             @I       J                 �Y8�?Z.��U� ?p             \@������������������������       ��;�4i?J            �R@������������������������       �%�;j� ?&             C@������������������������       �      d<             �?M       N                 `��?��}Qc�>k            �Z@������������������������       �                     �?O       R                 p�,p?S��'��>j            �Z@P       Q                 0/��?��|h��>             2@������������������������       ��.�O��>	             "@������������������������       ���#�)�>	             "@S       T                 �؉�?\��v��>X             V@������������������������       ��p6K�>E            @Q@������������������������       �h��2���>             3@�t�bh�hhK ��h��R�(KKUKK��h �B�  w+}��"?�j� Ec?�=Sj<�Z?�&����h�����)u��J#�ORo�?9�TN�&����_����d�݇��o�� ��g?U�I���u?5��g�?�PI���?�F�N$R?�n�;��׿�J���c�?�efd?Mܸ^��?��0�IIE��4�xp忽���z�?�����מ?Mm{?��?
TV���?\/����]?5Q�j�g?���!M}�17�H��?'0�ip#q��Y�����bO�
���?z����M�?��[���?@����?�X/ɢ��?+�~u{�?���F��?@�.��s?
)[C�t�?�9�T
i�?��
�ߕ<��0�'Ka� U�G����͔֔���?��>�n��� ��F���W���m�快�'���Dq��z�|�B  p�p���&��s�.��U�x{tc?C:=���z?O�.p�0�?�oˆV`̿hej45q`�mT9z������?�MEB�Xh��N��4�?FI5Ye� �o����?뀒���n�� iY(�⿞�BoBu׿��ڢ�F?��f�b?��/72^?��M�B[��3�����?M�<-��>�U��b?b��t��?�k��Y�����69��?���kGR�g�Th���&�g��JP�[��a��g���8T�|�'p��Vd�[�l��C�?���I[快��ͬj忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kqh�hhK ��h��R�(KKq��h��B�         :                 ��?K7bEn�#?�           �}@                        ��׹?O�q���$?"            r@                        ���?�	6�$?�             l@                        0�H�?	!yE;$?�             k@                        ��+�?0�7���#?�             c@                        �֧�?dU��G"?�            �b@������������������������       ������ ?�             b@������������������������       ����v'>?             @	       
                 t��A?�t $\�4?             @������������������������       � �i���?              @������������������������       �����C�>              @                        �q�3?f�H�ga#?A            @P@                        �bS?<�d��j!?'            �C@������������������������       ����x`}?             @������������������������       ���[�P?              @@                        ��?v?�?)ܼ�!?             :@������������������������       ���aC��
?
             $@������������������������       �v���#?             0@                         �Mm�?�@{R&d*?              @                         ��?�.)�l?             @                        `9F�?l��n
?             @������������������������       �                     �?������������������������       ��$(�L�>             @                         ��G? �2N���>              @������������������������       �                     �?������������������������       �      ��             �?������������������������       �                     �?       +                  �<�?���v#?A            @P@       $                 ��%t?1�S��@5?             1@       !                 ܬU?_H�*�"?             &@                         ���?`�?�VG'?             @������������������������       �`͉�g�?              @������������������������       ���hC
�>             @"       #                 �w?������>             @������������������������       �tT�@�d�>             @������������������������       ��CD�õ>              @%       (                 ��@}?�t}_��<?             @&       '                 �/?  �sz>e>              @������������������������       �                     �?������������������������       �       <             �?)       *                  /Ⱥ?���%�W ?             @������������������������       �                     �?������������������������       �H�Fߪ�>             @,       3                  �?nHLFo~?0             H@-       0                 �U��>Q��֡�?#            �A@.       /                 ����?�x+�p�>             0@������������������������       ��:��>             &@������������������������       �w��H�>             @1       2                 �f�V?���)�?             3@������������������������       ���}y�(?             @������������������������       �4�[�ľ>             (@4       7                 ����?P%o�?             *@5       6                 @ 
�?��W
�y?             @������������������������       �����v��>              @������������������������       ���14S�>              @8       9                 {�j?���jC%�>	             "@������������������������       �                     �?������������������������       �j�.��>              @;       Z                  ��?����__!?�            �f@<       K                 �<m�?`,: "?V            �U@=       D                 �1�?*W|~C.?'            �C@>       A                 �ۙ�?�/�H�?             3@?       @                 аs}?.��w�?             *@������������������������       � �}��
�>             @������������������������       �$�����>
             $@B       C                 �^7�?�v}�T?             @������������������������       ��S�}71�>             @������������������������       �R�5��>             @E       H                    �?>;s�2?             4@F       G                 0֥�?�����?
             $@������������������������       �                     �?������������������������       �`��ａ?	             "@I       J                 �ڡs?��A�?�7?
             $@������������������������       �8za7��.?             @������������������������       ���"B�?             @L       S                 0�?�?!��x��>/            �G@M       P                 �/��?��&,�?             *@N       O                  ����?�������>             @������������������������       �                     �?������������������������       ��Mp,���>             @Q       R                 @9��?�_
0�>	             "@������������������������       �x	b���>              @������������������������       �`R��e�>             @T       W                 h��1?�i�x[�>"             A@U       V                  ���?��>"��>             5@������������������������       ��Ȅ���>              @������������������������       ���\��>             *@X       Y                 ��b�?�=��ݢ�>             *@������������������������       ��m++0�>             @������������������������       ����o�ٸ>
             $@[       b                 p��?ڎ���?`             X@\       ]                 �$I�?�N�mV%?             @������������������������       �                     �?^       _                  �x��?j03��?             @������������������������       �                     �?`       a                 @�?����j�>              @������������������������       �                     �?������������������������       �      �             �?c       j                 `RZ�?��Ac|?\             W@d       g                 pZ9�?�G%�_ ?2             I@e       f                 ��s'?����]?             :@������������������������       �L#n:.�?             @������������������������       �s7T�?             4@h       i                 �B�?/�u�V ?             8@������������������������       �                     �?������������������������       �
�)!�l?             7@k       n                 � �?G����9?*             E@l       m                    �? w��]�>              @������������������������       �                     �?������������������������       �                     �?o       p                    �?���$?(             D@������������������������       �y�v�� ?"             A@������������������������       �ͧl��?             @�t�bh�hhK ��h��R�(KKqKK��h �B�  �H�Y7&��f7�HQ��/oL�0�(3+]�dF��"��a�3?��x�+#��I�Um:�?g_x��l�Y�?�mN�M �?�h���?KJP��h��K��:y����!�o�?�x�wf��9/8��[?t��C�ڿP}1���?؃j��D�?�12��~?��?��;]�u�fAQb��?�9�Q�1j�} M�"b忍~ӓk�	����0�?!���Po�*�������ٗi���LbT��3ͨo$�忦�*�¿�L�k?;������?�[�B�b�%����Е���b�ҙ�����/j�
���g����>����0�<��XG��_��w��t]�B�0���>�@��
�k�<a��F�u�?(;�/�g?���� �?,�ӣ�l�����M�{���s�����1p���a ���忆2Ѷ��Z���gv忻�?�_�ƨӵUT?��|��j?!�mC�?Y�>�Z�U?B�)�us?�/&-���l��T-��?	�X�<�x���7�����J��?������?N)N}w"v?������?�"�w��?x�Z��?x�'�o2�?�l�;�7�?9$��>�:�}�$p?N���jX�"cJoYi�?�X�Pk�].|%Dz?$E�0�ȿ$������?�� BY�a��yO+�gn��%r=F��N��_�`�j��|x7?򘧫�s�?'�Et�b�C�
��zC���u�<��� ,r��ij�^����$�[忤�5 �ӈ��]u���2����_� [v?� �)�\�WB&���a?��".��?HA $su��Z���x���5�fM��O���ݿq��a?�_*	!�?ÂF�c��?T&	���?
�	 �NO?���� ���WZ3b�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KGh�hhK ��h��R�(KKG��h��B�         0                 �)�?���
?�           �}@                          p��?�i[R
?�           �|@                        �v�?�k��p�	?�           �y@                        0��?�;*���?           0q@                         ڕ�?Ok��6�>�            �e@                         	Ù?����_�>�             e@������������������������       �>R��ť>�            `d@������������������������       ����s���>             @	       
                    �?|�vރ"�>             @������������������������       � �e�}!0>             @������������������������       � �ݢ	P>              @                        P0��?-�L�t*?e            @Y@������������������������       �                     �?                        P��?��ZE��?d             Y@������������������������       ��V����'?#            �A@������������������������       �nE5�?A            @P@                        ���?	"Ri�?�            �a@                        �Y&�?P��o�?             .@                        (GW�?'�v?             *@������������������������       ��&{B���>             (@������������������������       �       �             �?                       �o|?00|ؒ?              @������������������������       �                     �?������������������������       �       �             �?                        �ˤ?���f�A?}            @_@                        ਵ�?�kMWD?              @������������������������       �                     �?������������������������       �      �             �?                        P�!z? ����?{            �^@������������������������       �U���P��>             @������������������������       �z
��w?v            �]@        '                 8݀t?|hE� �?,             F@!       &                 PT�\?t���/�'?             @"       %                 ��ue?ʇݻߡX>             @#       $                ��D0!?`zCZF>              @������������������������       �                     �?������������������������       �       �             �?������������������������       �                     �?������������������������       �                     �?(       /                 �2*�?�I�� ?(             D@)       ,                 T�Y? EQ2:��>'            �C@*       +                 �r>�?�a��|��>             3@������������������������       �҂���_�>              @������������������������       ���?"F�>             &@-       .                 `�Q�?~z]s ?             4@������������������������       ��1;��^�>             @������������������������       ���6
���>             1@������������������������       �      <             �?1       2                 �Q�?�؞�>�?             *@������������������������       �                     �?3       <                 ����?��1;��>             (@4       7                 в��?($�N�b�>             @5       6                   .p�? p����>              @������������������������       �                     �?������������������������       �                     �?8       9                 �m�? ����2�>             @������������������������       �                     �?:       ;                 �/��?`eѷ|�>              @������������������������       �                     �?������������������������       �                     �?=       @                 �D�澘;�m���>             @>       ?                 0#��?�8w�X��>              @������������������������       �                     �?������������������������       �      �;             �?A       D                 ���?�O[��G�>             @B       C                 @q8�?�1h� ��>             @������������������������       �@_FsS>              @������������������������       �      X�             �?E       F                 �J��? ,����D>              @������������������������       �                     �?������������������������       �      ��             �?�t�bh�hhK ��h��R�(KKGKK��h �B8  ��B���>�0Ƹ�V��O��0��BK��J)?<{���E����՛9H���L^��E�f�f�3�Y^?7D_x�Y�?�~&��g�?��B�b[? ȯ
�?֭�dV?������?׈�S�:a�/��:�R�p�6��~u��َ[�g�k��5��Y�����?eE�甿�2Vtd��?\)�K��D�D6boE� %����?�@����?�̴�d�?�,GFY�L�6H☥.�?��M�~>ƿ��	�[?@��X��/�s��q,�lN���X��.��U��:�9$V�c%�ŪW��ݬ)���śr�e?�5��Uc?�JqJE$?$=��c��XV`/o�?����?r?~.�M��?q�P���?c�ȥ�?9[��_�l?v�RZ��?�6i��v_?ͅ���s? VTۘ�}?�����w�?��V��?UKs�R�i?-���p�?�.k��b?��U�]�?�W�3e�?`I�y�["� 4���d�1L���k���g�Y忸���I?���H2?a�B��X�?���ܰW� �^��@Y?�A:]�?+ʞ�L^�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kmh�hhK ��h��R�(KKm��h��B�         :                 @�C�?�}��R?�           �}@       !                 )DW?��a��?T           @u@                        ��]"?�7���?\             W@                         �\�?���r�	?H             R@                          ���?y�s�_
?             2@                        ���}?	ۇ���>             ,@������������������������       �"�S��>             &@������������������������       �Ɓ�G;n?             @	       
                 �P�?c��@�?             @������������������������       �`���`@�>              @������������������������       ��1A~l��>              @                          .p�?�d���?6             K@                        ț�q?�D�$�	?              @������������������������       �`�� &�>             @������������������������       �T����>             @                        ���p? �+6?.             G@������������������������       �kKh>"?             4@������������������������       �|*�)��>             :@                        P�C?��]'b�>             4@                        @F��3���>              @                        �@�?H�h���>             @������������������������       � *IY>             @������������������������       ��S���Je>             @                        ���o? �� pe>              @������������������������       �                     �?������������������������       �      �;             �?                        ����?��kO�>�>             (@                        xԠ?�x)e�z�>
             $@������������������������       �\�Zu�>             @������������������������       ��O*�W�>             @                         ��Tb?�?d����>              @������������������������       �                     �?������������������������       �                     �?"       +                  �6�?�ߎ���?�             o@#       *                 ����?��W?"             A@$       '                 ��O?6�u�ɱ�>!            �@@%       &                 𕖃?��gp�>              @������������������������       �T%�Y�>             @������������������������       �      �             �?(       )                 `T�g?a+,*��>             9@������������������������       ��]s���>              @������������������������       ����. ?             1@������������������������       �      8�             �?,       3                 �Q�?D6/g:��>�            �j@-       0                  �ڦ?��ae�r?M            @S@.       /                 �֧�?/	u$��?             9@������������������������       ���Pp��>             8@������������������������       �      �             �?1       2                 �*/�?ĵ �f ?4             J@������������������������       ���G�B%�>             :@������������������������       ����w�?             :@4       7                   ���?s�,�H��>�             a@5       6                  x�?���K"?              @������������������������       �x)��2?              @������������������������       ��G��
�>             @8       9                 0�,�?�vH+�>�             `@������������������������       ����!*��>              @������������������������       �q >AC�>            �_@;       R                 ;��?)l�~?�            �`@<       E                 a;�?�3}m?%            �B@=       D                 ���?F��WYB%?	             "@>       A                  ����?��k�3+?              @?       @                 �(�E?��=��>             @������������������������       �                     �?������������������������       ���^�>             @B       C                  `s�?�U��9�>             @������������������������       �                     �?������������������������       � �x`�E>              @������������������������       �      (<             �?F       M                 0	X�?��6�5��>             <@G       J                 P��?�\���>             *@H       I                 �p�?�kw�ͨ�>              @������������������������       �                     �?������������������������       �                     �?K       L                 �2*�?���8�>             &@������������������������       �����W�>
             $@������������������������       �      л             �?N       O                  $M�?�ެ���>             .@������������������������       �                     �?P       Q                   E(�?$�ĉc��>             ,@������������������������       �/A��a�>              @������������������������       �B�Rg�İ>             (@S       `                 P��?��@va?_            �W@T       Y                 P�)�?�m���0?'            �C@U       X                 @c��?�U��;�?	             "@V       W                 �c�}?@cr���>              @������������������������       ��G����>             @������������������������       �L[���>             @������������������������       �       <             �?Z       ]                 ���?g�fF?             >@[       \                  Ʒ�?��IF��>             ,@������������������������       �������>             &@������������������������       ����o?             @^       _                 ���H?�*W��)�>             0@������������������������       ���E��b?              @������������������������       ����s��l>              @a       h                  ��?=Z�n?8             L@b       e                  p<��?`)P�	?!            �@@c       d                 ����?���XϺ?              @������������������������       �                     �?������������������������       �      �;             �?f       g                  Z��?���$�?             ?@������������������������       ���#'���>             0@������������������������       �WG��E�?             .@i       j                 06y?��њ�>             7@������������������������       �                     �?k       l                  �E�?4��tJ��>             6@������������������������       �<ɐ��>             2@������������������������       �<\���>             @�t�bh�hhK ��h��R�(KKmKK��h �Bh  L��j�D�?s�n�8�]9�ב�N?�j@�"?�N�5�f�7���lXQ�����N�?�A�ۺ����+A�����n�1d���Y��@�Ϳ~���.>R?"��A�$z?��4ŧ��?VH�wah�? _b�/�)?8{Ӈ�Lοgr��&�?�p�8o? E���X?U�2���R?�ƺ�]�?Q[�R�Y�?�[�e?�a��e�?�_�2�b�?`��,�u?�g��<r?���'�w�?��JMf�?��Ӊ��?�ad���?K�����?����YL��N�o��/�͞�a��蜸Pz�8C�x忓-��?��m_I2�<I��������?��4Ҵ׿�Lt0�濎�1GFH:��L�kQ?�q��9�l?a��^���?�����?f���U#��I�Jֿ�1Z0 �?o�|t�S��(�F{���b��濾�}_�b�`���ӱL�q���b��?�!`�,�׿&>�\i2G?.=��W%j?Tg�α�?�G���t?�//z�5?/�:0���˄��?��	��v�?�u2LȨ�?:Yw���?H��2�?��|L�V?I���]�p?@�g�Fo�?"I�L��?�q����?L��d{e?=)�����?�K�`��?��nKN����6��I�/b��>��?��?��F�`�0h�c� 1�ז#��]�,���`�{��ׄ��q����R��%D�k�sĵ���Jݻ��6����]d?��k��5�?�E0��?��AT�g�j�6�s�f]���W����#�*K?Qʬ���c?���ߠ�?����2n�?gz`����?^
�?7"\?����ʁ�ND�?�N&xЩW����T��ɬC��P��di�?ӿ�
����忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kgh�hhK ��h��R�(KKg��h��B�         0                   �G�?�(^z��?�           �}@                        ,*�����1j�r?@             P@                        ?#�?w,�Gh?             7@                        p�N�?�7�u�?             4@                          ���?6U�=��?             ,@                         h��?�?����>             (@������������������������       ������>              @������������������������       � ީԚ��>             @	       
                ��Xv?�	�1�?              @������������������������       �                     �?������������������������       �      �             �?                        `��?��k�t	?             @������������������������       �                     �?                        ��jm?���9G#�>             @������������������������       �@$�R@�>              @������������������������       �4�-�$\�>             @                        PA��?v��F0?             @������������������������       �                     �?                         �G?�?n�d[(S�>              @������������������������       �                     �?������������������������       �      ��             �?       #                 �n�?!~���' ?)            �D@                         �X?��վ�[�>              @@                        `ϷP?0&�Ҁ��>             @������������������������       �                     �?                           �?�h����>              @������������������������       �                     �?������������������������       �                     �?                         0?+HW8�h�>             =@                        P�c�?EtD�H�>             @������������������������       ������>             @������������������������       �                     �?!       "                 �ڡ3?���_՚�>             7@������������������������       �                     �?������������������������       ��"+�q�>             6@$       )                 ����?��i��	?	             "@%       (                 p۶�?���q�>             @&       '                 �_��? �İR�>              @������������������������       �                     �?������������������������       �      �;             �?������������������������       �      �;             �?*       -                 pM�T?��T��>             @+       ,                  �Q�? '���qy>              @������������������������       �                     �?������������������������       �                     �?.       /                 0n�W?_J��>             @������������������������       �                     �?������������������������       ��{2��z>             @1       J                  ����?�z�Jl?�           �y@2       ;                 `f��>ʃ}9 x?�            �k@3       8                 ��`�?�"�Э�>             @4       7                  �vg?P$A����>             @5       6                 @F����WV�>              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?9       :                 0�!�?���~�F>              @������������������������       �                     �?������������������������       �      x�             �?<       C                 �\ͥ?��C[f?�            @k@=       @                 ~`��^�	�R��>             (@>       ?                 ���?@������>             @������������������������       � �%M �>             @������������������������       �                     �?A       B                 `��?�+�DX��>              @������������������������       ��W��m�>             @������������������������       �      �;             �?D       G                 @Ws�?�l/L(�?�            �i@E       F                 ����?�*A�?              @@������������������������       ��QS���>             .@������������������������       �Lx�;�?             1@H       I                 �k��?L��SB?�            �e@������������������������       ��\�{��?             @������������������������       ���|�R?�            @e@K       Z                  ��?Q꓉<?�             g@L       S                 �Lj?�.���?~            �_@M       P                 �xb?�R�s�2?             *@N       O                 ���d?��$|��>
             $@������������������������       ��-;�8P�>              @������������������������       �X��VЙ�>              @Q       R                 g�a?`�V���>             @������������������������       �`a��J�>              @������������������������       �      �;             �?T       W                 𤔭?Z@�X?q            @\@U       V                 ����?2���K?*             E@������������������������       �kwaDh>?%            �B@������������������������       �7�k�2
?             @X       Y                 �C`�?
�عk?G            �Q@������������������������       �T���C�>              @������������������������       ��se��<?E            @Q@[       `                 �o�?�;��M?;            �M@\       _                 ���?���
XL?             @]       ^                 ���|?<��M\��>              @������������������������       �                     �?������������������������       �      ��             �?������������������������       �                     �?a       d                 @J�?��ҥ?8             L@b       c                 �\��?h����
?             <@������������������������       ��J�He?             9@������������������������       �D�pr~?             @e       f                 @� ?����|�>             <@������������������������       ��|��
?              @������������������������       �BN�pgq�>             :@�t�bh�hhK ��h��R�(KKgKK��h �B8  �C���k	?[bwY?�/���s?�K.A�;f?'�{۵r?I��g?oIr����?�<Ǚ~�?��%��ߍ?���IZ��?u��i��?WS��fZ������(Kviq�S?�#�,Ed�h��Mm�?5\�Rq�?�*�=4�?@����"{?vg����?� ~!b�?�>�SBy,�R�J�/�F?
���Z�s��,v^�X�?�^qBq�~�d 8�A�心��<jw忬�Ώ��T?�^+Üe��F+�_����r��q�%J��b?�@Pl��?<c׻���?��ҙ[-l�X��'����Ղ6�q��0����0 ."܂�7a-#������,O?����@l?�����f�?��	`�i�?�ha�{3���mdeY�?��I��Y�b��j(��&���H���T]�dr?+���4�?�8���
z?�k�kt�?4��#|�?װ��5��?���q1E�O���HX忹�KjY��d��K�;,A1q������������!@���*�Kp忎%��'@\��D>)m��O��y�?��T��E���5w_�Y? ���WԿ�n�k_�?�����Q��AH#���\-Џq��i6ҁ�\??[�= �4�"�0��m?��m���B?*A��Ŀ�z���t�?U��3 #�?�`)��?i�((�|�?0���?I����sfd��n�PCۿ��ޣ�?)�\A,0?��'��?@/
Ð�;�c�'�a?�k����?RFg�r�X�a���U忤��d�e���X���?�Ĭ��T?`;�Xl?[�m�d�?Ӣ���?Y@�)!�L�HK��U�?��#i`࿔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K;h�hhK ��h��R�(KK;��h��B�         0                 ���?&��@�>�           �}@                         Z��?B5��S��>�            }@                        `TF�?4k]����>�            {@                        @E��?_�G���>�           {@                        ��P�?��Hƍ�>K           �t@                        ���?��=�nX�>4           @s@������������������������       �[���qW�>/           �r@������������������������       ��筩?             @	       
                 0Ղ�?O�]go�>             7@������������������������       �                     �?������������������������       ��ت��|�>             6@                        `RZ�?� T8P�>f            �Y@                        �#;�?##��}��>             ;@������������������������       �hz<��/?             @������������������������       ����뭖�>             8@                        ���?���ꒄ�>K            �R@������������������������       ��û�n��>	             "@������������������������       ��m��Z0�>B            �P@������������������������       �     @T�             �?       !                 `�??�N�7�>              @@                        �Cl?��+�#�>             6@                        �Ƹ?9gF*�>             0@                         ��e?"�+ǉ�>             ,@������������������������       �8%)�S��>             @������������������������       ��D*�B�>	             "@                         �a�?D��%�ְ>              @������������������������       �                     �?������������������������       �      �;             �?                        P�~x?��rA�>             @������������������������       �                     �?                          ��?�)%{Tc�>             @������������������������       �p�L	d�>             @������������������������       �vذ�wv>              @"       )                 �dŀ?X��E� ?
             $@#       &                 h��?�q���'�>             @$       %                  ��^�?@��~=�>             @������������������������       �                     �?������������������������       �  �Ru�W>              @'       (                    �? �G%��x>              @������������������������       �                     �?������������������������       �      �;             �?*       -                 в��?�B��_��>             @+       ,                    �? A(��N>>             @������������������������       �                     �?������������������������       � x��g�">              @.       /                 ���?�+�����>              @������������������������       �                     �?������������������������       �      X;             �?1       2                 ���?�eG��>             @������������������������       �                     �?3       4                 p��?�c4"\�>             @������������������������       �                     �?5       8                 �P��?'�@�`�>             @6       7                   ���?����>              @������������������������       �                     �?������������������������       �      P;             �?9       :                 ġl�?Ζ �Xh�>              @������������������������       �                     �?������������������������       �      C;             �?�t�bh�hhK ��h��R�(KK;KK��h �B�  �&�:�>ۗ���(��Z �?��}���?���r
)��к�;�
����m 1�?^��F��࿖�}'<�`��0u����"�Q>Bݿ�:�48 J?,��a��c?�H�09�?Ӿ�`r�?o���KG,?������m-�j�?j"��|��?�r��B�W����-)����LeFJ�;�ب�T���qh��ɿF�*a忀H^�N�a? �Oɬ[�?B�5�f�?�ٞ5:~W?�8k�7e�?f|�AC�R?իAY�^�?Ic�X�?��(�vCq���x�y����"ͯ��lۆ�(��y�+���lF��uh��Y[g忒Q� �c忓Q��? ��	_R?�7��
\�?�0ǡ/[�?A�S��RW���kC\f��-[�V�?\��yվk?�aH�I��?�j�	OS?&���n�?T��~C4? eI�F�Q?����]�?K��X�?X���>����F�Z�C��U�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K7h�hhK ��h��R�(KK7��h��B         6                  @���?D�s"�L�>�           �}@                        �x�y?^�����>�           p}@                        ����?h��ޒ}�>	           �p@                        0�?�?CJSq��>�            `d@                        ����?{v� m]�>�            �b@                        �=E?�F-�q��>�            `a@������������������������       �"k9�|��>o            �[@������������������������       �tf6��>             <@	       
                 �u�?,@����>             (@������������������������       �                     �?������������������������       �> �����>             &@                           �?��1^�?             (@                        �o�?��mX$�?             @������������������������       ��{��>             @������������������������       �`�����>              @                        ��ى?�n�1O�>             @������������������������       �  �K��=              @������������������������       �2�f=���>             @                        � D�?��s��>f            �Y@                        P���?i���E�>:             M@                         �\�?��/��6�>9            �L@������������������������       �&{	�(��>             &@������������������������       ����>�>.             G@������������������������       �      <             �?                         �g<�?Z�kR���>,             F@                        `@��?� �A/�>
             $@������������������������       �h�i�@��>             @������������������������       ���e^>             @                         a�? ?����>"             A@������������������������       ���b��Ȝ>	             "@������������������������       ��&��t>             9@        -                 �D�澽~���M�>�            �i@!       &                 ���?mS�պ ?<             N@"       %                  �Ѱ?l�B� ?3            �I@#       $                 �v��?�NȖaR�>2             I@������������������������       ��5���>'            �C@������������������������       ��4�����>             &@������������������������       �                     �?'       *                 ���?�����>	             "@(       )                 ����?�� Nܛ�>             @������������������������       � �f�)j>              @������������������������       ��t͉��3>              @+       ,                 ��?�?ة��7�>             @������������������������       � �8y�k>             @������������������������       ��@�cP�>              @.       /                 �z?�P�-׬�>�            @b@������������������������       �                     �?0       3                  `s�?�����>�             b@1       2                  �6�?K�$��>             @������������������������       ����12�>             @������������������������       ���
?��>              @4       5                 ਮ�?����-�>�            �a@������������������������       �3�c�dl�>3            �I@������������������������       �؋�(���>Y            @V@������������������������       �      /�             �?�t�bh�hhK ��h��R�(KK7KK��h �B�  �x?�6�+q^Z��;����>��C�"��x��6�6���0᩠$�_�K��D�?�2����׿���.��d�+ �������ֿ;>���c?��?Ѥ�t?�����?N\�x���?� ��OHU��/�{�k�|��C�?4�}DjXP��c�kݱZ�V"R�\X��S5�r�?Н�b����������_��%��Z�F?�}k�j�?1��"�W�T��]�];�g7�]�w��nuX���p��7?�-��/^?.�J�X�e?��"�`?&*\ޔP�?�7�d�t��Fu�?��s�?�f��ħ=H�� l��\忸v�YV忔;��q�p*4f�g�"ׇz忲��Y�00�1^����?i���5�Z����Ef?��n}K�?y���u�?Y2����<��]�
{�׿O�e�ǚ��~j�Y��?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KOh�hhK ��h��R�(KKO��h��BH         2                 �jx?s愎���>�           �}@                        @j��?�5K��V�>           �p@                        0�I�?I�4�$8�>�            @j@                           �?R��>��>�             j@                        p�t?D���;��>�             a@                         .s�?�*�#��>�            �`@������������������������       ��A?��T�>p             \@������������������������       ��;a�p�>             6@	       
                  �a�?���N�>             @������������������������       �                     �?������������������������       ��Hj	�>              @                         ��^�?N��J�>G            �Q@                         y��?�O~R���>5            �J@������������������������       ��]�	�"�>             1@������������������������       ��f��b��>$             B@                        �j��?J.eL�~�>             2@������������������������       �.}��b�>             (@������������������������       ��� ��O�>             @                        �۰�?���^H�>              @������������������������       �                     �?������������������������       �      �;             �?       #                 ���?��d��|�>6             K@                        0?��Z�7�>             (@                        �@�?`^��:�>              @                        0�,�?�b�|���>             @������������������������       �                     �?������������������������       � ��O4]>             @                        �@I�?`�u�0Q�>             @������������������������       �pfh�4�>              @������������������������       �   ��x=              @       "                 @��?̱�(A�>             @        !                 0׆�?@@ZjP>             @������������������������       �                     �?������������������������       �  ԡ]Ek=              @������������������������       �                     �?$       +                    �?[��
���>*             E@%       (                 �ζ�?��l�_�>             .@&       '                 ��M�?Ї�J�>              @������������������������       �                     �?������������������������       �      �;             �?)       *                  p�Z?����t��>             *@������������������������       �V���j��>             @������������������������       �|��%9ǝ>             @,       /                 ��?�2��f��>             ;@-       .                  �Mm�?j(>�L��>             @������������������������       ��p)�f��>             @������������������������       �@�X���O>              @0       1                  ���?5g�7�f�>             6@������������������������       ��+�`��>             (@������������������������       �
?H/|��>
             $@3       8                 �z?��vJ��>�             j@4       7                 �T�?��_��>             @5       6                 �d?@�i�F��>              @������������������������       �                     �?������������������������       �      �             �?������������������������       �     �Ի             �?9       B                 ���?�xH�g�>�            �i@:       A                 ��ذ?j5���x�>�            �a@;       >                  �8�?�w�IbG�>�            �a@<       =                 `��?]�(��]�>�             a@������������������������       ��y�i�>              @������������������������       ����XW�>�             `@?       @                 pp�?V�Ph~��>             @������������������������       �L���ϕ�>             @������������������������       ���ж�	�>              @������������������������       �      4�             �?C       H                  ��?O���P�>>             O@D       G                 ��L�?��:B��?             @E       F                 `۶�?�:f�p�>              @������������������������       �                     �?������������������������       �      ��             �?������������������������       �                     �?I       L                 �D��b=�7��>;            �M@J       K                 p���?X� �>1�>              @������������������������       �<$s81�>             @������������������������       ���Q��;>             @M       N                 ���G?�q���f�>3            �I@������������������������       ���YةC�>             @������������������������       �Rv
W�B�>0             H@�t�bh�hhK ��h��R�(KKOKK��h �Bx  "M�F�?��Z'�<?�I`x9H?W�l���E?4�oF�,?�V[v� ?rA�YV��?��g�#Sӿ+��9�q?P��b�?���k�q�?��<�X?�f5�a�J?��t�M�ο��ֵ�?��� m?ǤB2��?F�CL�?@��:2�?�Fc]f��?.KY�9��?�
� �G�U�7�8`g���<��n���}���s���O�vk�&���q�$l@�7e���q�U_��+�'h�>#Oi�6R�e��4�W4��<A�V�1�MāW����h�ZQ�ЖR�@@���\^? Z:��5�?�]<[ߘ�?���~�?ETt�RD?FO�#�?*���o]忛��g��S��e�R�q�߭~h|�����Z忢1��{@�"�U����?���M���}����8�cR4��{���U�B��� g�E?�忀�v����hW��T�'�2�'+��%G� �$nTf@�/��D��|3*��?���Z��ȿ�
���k?INP{Z�g���X��?� �����
MndF?U¨��|? �X��d?���9�h�?<Q��a]�?>��l9��?��l8��6?�DY)��m?�ۏ�r��?Ĥ(��Y�f@{&�r%����dw�$=�,�x�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K#h�hhK ��h��R�(KK#��h��B�         "                  @���?�J?�%��>�           �}@                        ��g?���2Z�>�           p}@                        p4 �?�U�cV$�>i           �v@                        �)�?"d���l�>h           �v@                        ���j?p��V[$�>`            v@                        0�B�?x������>�            �l@������������������������       ���-���>�            �h@������������������������       ����{;��>              @@	       
                 0]��?���A�>y            @^@������������������������       �G&W�V�>w            �]@������������������������       ���i���>              @                        4 �?�:�i\�>              @                         h��? �%�s�:>              @������������������������       �                     �?������������������������       �      ��             �?                         X3�?֭�^��>             @������������������������       �P�k�Ń{>             @������������������������       �x��'c|�>             @������������������������       �     �0<             �?                        ��I?�4����>n            �[@                        pS�j?g�� ��?              @������������������������       �                     �?������������������������       �                     �?                        Ў m?\_�K���>l             [@                           �?@����?             @                        |ِ?�e�
x>              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                        p�m?�_C�V��>i            @Z@������������������������       �                     �?        !                 pJ�q?�f���>h             Z@������������������������       ��`�܏��>             @������������������������       ��<��>c            �X@������������������������       �      �             �?�t�bh�hhK ��h��R�(KK#KK��h �B  d]�h��e.9�\�>��K5z�&�u�2�)��g��s/���t�C̾.�|��Z��?k�#/�?$>Vb7�F��` �s�Ϳg�ٔ��5"���[?@.�K`�x?7V1��u�?�I�p�v�?q*� B2?�H�8Y�u����\�?p��s��?ّ�1�D? �5��a~?�]4r[�?�4I��?�;$�@?�bȩ�f� �k���V?��c�_�?{��Z�?�ʗ�C���y$���C?F]iGw��?�B;�T@?l�=�KP࿼����?�Z�WA�忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K3h�hhK ��h��R�(KK3��h��B(                          @I�>jN����>�           �}@                         `���?������>             @������������������������       �                     �?                        QU�>$ژ"xտ>              @������������������������       �                     �?������������������������       �      ��             �?                        �߯�>r�]@֌�>�           P}@                        ��xg?"�<6I�>             2@	                         �ǽ>q�\�*�>             @
                        0� ?�w���>             @                         ��>`+�-�>              @������������������������       �                     �?������������������������       �                     �?������������������������       �      ��             �?                         ��d�?�(��m��>              @������������������������       �                     �?������������������������       �                     �?                        ��'|?�1�����>             *@                        �m�?��&j�۸>             @������������������������       �                     �?                        �T?`����Kv>             @������������������������       �                     �?������������������������       �  �6��=              @                        �m۶?�c���s�>	             "@                        ��?ƽ��'-�>              @������������������������       ��xF[�߿>             @������������������������       �����_�>             @������������������������       �      »             �?       $                 �D�>l�J��>�           0|@       !                  `���?�d�?             @                         _5?ܼ�l�>              @������������������������       �                     �?������������������������       �                     �?"       #                  `���?[`4���>              @������������������������       �                     �?������������������������       �      ��             �?%       ,                  ���?�m�6z�>�           �{@&       )                 P���>�ۂ��>!           r@'       (                 ���q?�i�?9Q�>              @������������������������       ��@TR�ʸ>             @������������������������       ����k6>             @*       +                 �"��?*����>           �q@������������������������       �� pp3��>�            �e@������������������������       �ϴѶ��>l             [@-       0                 `�Q�?�{��Y�>�            �c@.       /                 ���?
ãG��>*             E@������������������������       �{�w���>(             D@������������������������       �@�%H��>              @1       2                  @���?2?ԁ*�>t             ]@������������������������       ��Lƪ+G�>s            �\@������������������������       �      �;             �?�t�bh�hhK ��h��R�(KK3KK��h �B�  id᭗�> g}Մ�o?��
{�?���L0�c?��R��i�?��f��Z�?�e��C��ب#R��Z(r��:Eh�T��j|���f�^�4Yh�ɣ)�`����_�?�:{.����|/!Ǘ�f�o�w�'�J'�h&? `��Xn`?�I|ӥk�?UG���U?����^�?�y�l[�?j��rAE�,���2�P�6/:�d�>(L>�~�?�@�b�?�a;��i�>rC��FMk?8K�B:^�lmЖ]�?0
�g�q� �.�jg�?�c��T��?����q�?\ArB��>!4ӆ�e'?a#�/�_�V`��i忹�C�~W�?��+�B/?�����b�?�=�{&���5j��R5��q��O��f��]Ŀc�Ɏɑ忟�=/�٠PJ��ƿ��k��l�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K?h�hhK ��h��R�(KK?��h��B�                          @I�>�/��8k�>�           �}@                        �y���^���}�>             @������������������������       �                     �?                        @1e?p��^��>              @������������������������       �                     �?������������������������       �      �;             �?                         �C[?�GѫL�>�           P}@                        pF�T?�@�L��>             >@	                        �/��?�^A{���>             ,@
                        ��IL?��UTH�>             (@                        �h�J?�݇����>             @������������������������       ��^V��۬>              @������������������������       �      �;             �?                        ����?p�oƠS�>	             "@������������������������       �0���^��>             @������������������������       ��g#<g�>             @                        `��?*��1���>              @������������������������       �                     �?������������������������       �      l�             �?                          .p�?�t���>             0@                        0�?5=�kiN�>	             "@                        (�&R?�O�q�S�>              @������������������������       �                     �?������������������������       �      �;             �?                        @Ws�?��7��>             @������������������������       ���Xԍ�>             @������������������������       �@&Pv2=�>              @                        x�8a?��uj��>             @������������������������       �                     �?                        ��eS?���"�/�>             @������������������������       ���囇>             @������������������������       �      ��             �?!       0                 ��Zy?�\$�>�           p{@"       )                 �0l?ɕ7f�^�>K            �R@#       &                 x�S?��9��>,             F@$       %                  ��m?��0$��>              @@������������������������       ��O�.���>             3@������������������������       �%,1̒��>             *@'       (                   +Y�?z���5s�>             (@������������������������       �??)�>             &@������������������������       �      �             �?*       -                 PQ�p?0N꒛��>             ?@+       ,                  P��?0�$��>             @������������������������       �                     �?������������������������       ����`��>              @.       /                 �><r?�;Ԃ�g�>             <@������������������������       �                     �?������������������������       ���I�;7�>             ;@1       8                 `��?i�Ń8��>l           �v@2       5                 `��m?�f�S��>1            �H@3       4                 �x�?���Ǳ��>             8@������������������������       �� �S��>             0@������������������������       ��-N�=�>              @6       7                 `�?��g6���>             9@������������������������       ��~����>             8@������������������������       �      �;             �?9       <                 �c��?�\�F���>;           �s@:       ;                   E(�?�u�ߵ�>	             "@������������������������       ��O8��/�>             @������������������������       ��\��>             @=       >                 *��>���Y��>2            s@������������������������       ���=$��>              @������������������������       �Jta|���>*           �r@�t�bh�hhK ��h��R�(KK?KK��h �B�  }&h]��>ŷ��No���pYz忋�<z�bc����i��K��Z�)��l��>\����R?~�{X��d?|Z(�*�i?����MP?�ůkh�?3Y�6h�U�4���o?�Լd�s�?0���7e�?���*�U��;hѼa�ϳ�tW�j)��1�#�GfZ�~JY���{�[u�K�8����(<:�gc�r2;k7@�l<�u���?Q�XKj�SiSK�Z?G�l�p^�+��[�a?�_�?Cb�#�l�?�;Ğ���D�F~+E����vRV��br0+;����H��?Y`��y��>��o��ޢ�t�;�j�快�vUL8? "N�rn?YB�!�Z�?]~�lq�?ɩRB���>��@|�,a6��8�?<�7
�?0ri oR?Gi��_?y��Sh�?��J�t�?��<��2?��1r� m�p��*3~�?&�p�����v���d�.��C��忝�fE�?�Sg�_ܾQƿ���T>��A�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K_h�hhK ��h��R�(KK_��h��B�         0                   s��?N �/;�>�           �}@                        pҷ?�ʭ����>�            �e@                        ��e�?�/#[v�>w            �]@                         ���? �8�IӠ>o            �[@                         '�?��TUr�>n            �[@                        P��?�x�W9�>k            �Z@������������������������       �t62u���>e            @Y@������������������������       �쬂�Gj�>             @	       
                 �'U�?�\qd��>             @������������������������       �'ض�Kc�>              @������������������������       �      ��             �?������������������������       �      ��             �?                        ��A�?F�{���>              @������������������������       �                     �?                        0vb�?��:/K�>             @                        �2OF?"�KP֗>             @������������������������       ��)̾�r>             @������������������������       �                     �?                        �x��?���鋷>             @������������������������       �@a6(���>              @������������������������       �      ��             �?       #                 Px��?$�L�29�>8             L@                         ���?�L�����>             @                        P��;?�f�C��>             @                        ����? ��qoM>              @������������������������       �                     �?������������������������       �      �;             �?                        0��?�[�;41)>              @������������������������       �                     �?������������������������       �      P�             �?                           E(�?���QÔ>             @������������������������       �                     �?!       "                pT�? <lD�p>              @������������������������       �                     �?������������������������       �                     �?$       )                  ���?t�� ��>1            �H@%       (                 ���?�<j��>             8@&       '                 pM�D?�HV����>             7@������������������������       �@�Fuq�>             *@������������������������       ���[v��>
             $@������������������������       �      �;             �?*       -                  ^ߵ?NoҜ=�>             9@+       ,                  �9��? �����=              @������������������������       �                     �?������������������������       �                     �?.       /                 pD�?�i���ı>             7@������������������������       �Ɛ�4�>              @������������������������       �~k����>             5@1       B                 `s5�?SV ���>)           �r@2       ;                 `Fe�?I�a�/�>             ;@3       :                 𱯬?����)�>             5@4       7                  ���?}�S� Y�>             4@5       6                 Ȇ�d?�~��c>             2@������������������������       ����5�\>             0@������������������������       �������>              @8       9                   ��?�1�S��>              @������������������������       �                     �?������������������������       �      �;             �?������������������������       �      �;             �?<       =                 p�_r?�IC�2p ?             @������������������������       �                     �?>       ?                 �\ͥ?� ����>             @������������������������       �                     �?@       A                    �?�W!�iQ�>             @������������������������       � `�����=              @������������������������       �����z�>              @C       R                  /Ⱥ?�p�]Xv�>           �p@D       K                 ���?���63{�>x             ^@E       H                  ��M�?�C��>n            �[@F       G                   �g�?���O�!�>i            @Z@������������������������       ��}�Q�>g            �Y@������������������������       ��!D�u��>              @I       J                 (OUC?D[QT��>             @������������������������       �gRJ���X>             @������������������������       �                     �?L       O                 ����?�����>
             $@M       N                 0~��?�&���>              @������������������������       �                     �?������������������������       �      л             �?P       Q                 ��d?�EV�}�>              @������������������������       � `{��|[>              @������������������������       �hy/훐>             @S       X                 pk�?ب�����>�            �b@T       W                 �nN�?��U�mb�>,             F@U       V                  �~��?x6g3��>+            �E@������������������������       ����P?              @������������������������       ��o�A�>)            �D@������������������������       �      �             �?Y       \                  9ר?�á�Y�>j            �Z@Z       [                P�ᨪ?�Iߙ̄�>              @������������������������       �                     �?������������������������       �                     �?]       ^                 @��8?G��	�>h             Z@������������������������       ��&�̽
�>$             B@������������������������       ����V$.�>D             Q@�t�bh�hhK ��h��R�(KK_KK��h �B�  +��J���Ʌ��{1���P �"��� p�-�G��	I(��`.x�c-��L��n�ݿ�65�%^忣j
�*�S?V,�y���?�m7�/c�?��H�Oo�v��+?{b?� ؔ��?�F��{>?R8fbHL�GT{�X�՞�_I_� �i��2b?Ǔqcf�?��MKY�?�N��	/G�x$?t��d�K�``��H��cGJP�S��$'�\�e#0�7[忺BfX�5�� !�V�o<��bW�+׎w� t�!��l�s�	�o�u��̙�s�`�`��p�{A�nX=�Y���}�Q�@]v�N�ݜ���c�9e�9�=տ;��h�m�����$?��[�,c?�m�Db�?_�Ȍ,b�?�6�g�d��u�D�(h�?t�..^Ͽo1<G�G!?z��v"�L?4/�Q7� ��2����#?�r�{��p;�O&W�2�҉V�? `�u�c?{yJ��l�?����TX�?�J�i�E染p?��"r���?-�f��5]?����Dz�?���*�A?|�AP]�?�QS�ܿ�M0?�	���0���Y)��C	
%����Ŀ�lp�+��{�AS?F�~��V忩S��x�?n��,.<^��i�v����*.g�{#���|�u8;�M��R%;bd��8PV�ڿ�r�ب�3?���[S?�荿pO?����J�?��j����?o�W	���?m���rK��+50��w��ؐ�`忘^�f���N�a�?_������?|���Wd���t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KQh�hhK ��h��R�(KKQ��h��B�         6                 @�C�?Y���L<�>�           �}@       !                 ���u?�/ld��>T           @u@                        p'v�?b��}���>�            `a@                        �U���F�v~��>s            �\@                         ʟ�?�銬6�>1            �H@                          ��?d������>             3@������������������������       �=]c��D�>             1@������������������������       ���_j͌>              @	       
                 �J ?}��Н��>             >@������������������������       ���O�à>              @������������������������       ��F$�i��>             <@                          �x�?�9��>B            �P@                        P+�Q?��y)���>*             E@������������������������       ��4��h�>              @������������������������       �����2�>(             D@                        `Fe�?+����ܻ>             8@������������������������       ���c4!��>             *@������������������������       �9�z��>             &@                        `�X2?&D��D�>             8@                        `焘?޻Z�2J�>             *@                         `�J�?��Я��>
             $@������������������������       ��|�俢�>             @������������������������       �������>             @                        �qht?�F��ꬪ>             @������������������������       �  ��R0>              @������������������������       �      ��             �?                        ��,P?y]���&�>             &@                        ��T<?~��z��>             @������������������������       ��A����>             @������������������������       � c)�P6�>              @                          �a�?�*��F��>             @������������������������       �Z/�ҵz>             @������������������������       ��|=�Or�>             @"       +                 �Z��?7`��7Y�>�             i@#       *                 `���?|���\�>&             C@$       '                 �I?�*�U���>%            �B@%       &                 �p�?�_�����>             6@������������������������       �ʕ��?1�>             1@������������������������       ��~��Ff�>             @(       )                 ��>}?ePR�>             .@������������������������       ��;TGI��>             @������������������������       ���]<��>             (@������������������������       �      �;             �?,       /                 p���?V��?�>�            `d@-       .                    �?� ����>              @������������������������       �                     �?������������������������       �      ��             �?0       3                 �{��?��A����>�             d@1       2                 0��}?�MHf��>h             Z@������������������������       �Bj�ӣ{�>             &@������������������������       �3E�Xj��>]            @W@4       5                   �P�?Q5/����>9            �L@������������������������       ��96�%�>             5@������������������������       �z��o?�>$             B@7       8                 ��r<?�l#hy�>�            �`@������������������������       �                     �?9       B                 p��?�3s����>�            ``@:       A                 0�0�?�&T
b�>)            �D@;       >                  �^�?��v�1�>(             D@<       =                 *]�?����a�>             ,@������������������������       �����Ҽ�>             @������������������������       �nȔs��>              @?       @                  iB�?��M��>             :@������������������������       �ؾ�����>             .@������������������������       �v[�IE5�>             &@������������������������       �      �             �?C       J                 `WJ�?+��u(I�>Z            �V@D       G                 ����?�kɕ���>1            �H@E       F                 `�Y�?�۱�欭>/            �G@������������������������       �,)t� ۪>             >@������������������������       �V�Ѝi�>             1@H       I                 h��Q?g d�z�>              @������������������������       �                     �?������������������������       �     ���             �?K       N                  ���?�������>)            �D@L       M                 �'��?Q�D[�>             @������������������������       ��IpA��>              @������������������������       �                     �?O       P                 �Y8�?�r|s�>&             C@������������������������       ��\�W8�>              @������������������������       ��(���5�>             >@�t�b��      h�hhK ��h��R�(KKQKK��h �B�  io(�ˆ�>v��7��\��!6�$?ŞB>�K��(�d�3�E�1�����:?�6�)��?s���b��M� KV��o��p�b�F,�ٿD#�t�=?��K|�!?�h~Hd�K���w�?_at'}�P?�T�[&��?TR����?�TM�P?� a�`?�L��T?0�V�_�?t6��Z�?�!�"is?��k�r�?y�gh�?S����)��J1��bU����2�?���dh�OX��G?�	��X忊�FV���?� ����0�ㄗ��P��I���H���[��9^�@�>���п�SE�z�������K?�Cƥ�n�?�k��;�?�ѫ�Ԏ�ě|�!�@��)up?g�u�Tg�?�#T�go�?�{���!����_7��G �`�H�Eŭ�ӿ�/	a.�1?V�ޑ�;�?��j&/�ƿ�ڮL�5?�UJڢo��
sc�{8?� ,�
�P?>�>�@�M?%=,@Q�1��ER��?7Ħ ۿp�L-�W?I��,f�?d��>��?"���v�?������?�R�hq5��5��-�0�H�ŕ޿!�B`�?[kC���e��I5/r�e��s�U��Kn�n�A?����s?C�7J�@�?�C;���?�u��O,?J�-q���?Mm���KϿ�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kwh�hhK ��h��R�(KKw��h��B         :                   s��?��Tb��>�           �}@                        ��a,?�Έ�(��>�            �e@                        `q��?$U:�*$�>\             W@                        �w�m?g�����>7            �K@                        ��IL?�<=d��>             2@                        X��?2\����>             @������������������������       �                     �?������������������������       ��Q�;u�>             @	       
                 (	2?������>             ,@������������������������       ���9��>             @������������������������       ���f��B�>              @                        ��N�?��oLO/�>%            �B@                        �$I�?��9�h��>$             B@������������������������       ��=<�#�>#            �A@������������������������       �      �;             �?������������������������       �      ̻             �?                        ����?s�L��>%            �B@                        �p�?Pi2�&��>             @                        @"��? ��Z�9�>             @������������������������       �                     �?������������������������       � ����P|>             @������������������������       �      ��             �?                         ��g�?��%���>             ?@                        0���?O��vY��>             @������������������������       �8G��ߵ>              @������������������������       �l��;���>              @                        0}}?J��u��>             ;@������������������������       �>]j7��>             @������������������������       �QU1�A��>             8@       -                  �\�?�`ii׊�>S            �T@       &                  G8W?�Ӣ�V�>*             E@        #                 ;��?y��F��>             @!       "                 � �?��i�z>             @������������������������       �                     �?������������������������       � g#��5I>              @$       %                  �0��?��O��h�>              @������������������������       �                     �?������������������������       �                     �?'       *                  ��i?ۤ����>%            �B@(       )                 �۫e?@z?g��>             @������������������������       ��-� B�>              @������������������������       �                     �?+       ,                 �>��?��`OJ�>"             A@������������������������       �~�$�;�>             6@������������������������       ��{7֠�>             (@.       5                 `��r?�*��e�>)            �D@/       2                    �?��Ӎ��>             ?@0       1                 �@�?`C�!;�>             *@������������������������       �,ѩ_�>             @������������������������       �l�&�*k�>             @3       4                 (��@?�-^B��>             2@������������������������       ��օ�R�>              @������������������������       ����)�>
             $@6       7                   ��?��v��>
             $@������������������������       �                     �?8       9                  6��??7y}��>	             "@������������������������       �Zž��^T>             @������������������������       ���Ǭ�Q�>             @;       X                  ����?7����0�>)           �r@<       K                  �/�?�_P���>p             \@=       D                 �؉�?�ɫ�!��>&             C@>       A                  m�a?$���7:�>             0@?       @                 HR	 ?��Y@p�>             @������������������������       ��z�R��>             @������������������������       �                     �?B       C                 ���@?�#V��>             (@������������������������       �0�kOd��>             @������������������������       �ږSF�>             @E       H                  ���?�Q��_��>             6@F       G                 `U�?�<y����>             .@������������������������       �`�y���>             @������������������������       �H��r���>	             "@I       J                 ����>���JY�>             @������������������������       �                     �?������������������������       �}���
�>             @L       Q                 ���?��	.���>J            �R@M       P                 �ǔ?L��;�+�>             ?@N       O                 \F�M?@�{�>             >@������������������������       ��i�KP�>
             $@������������������������       ���pyX�>             4@������������������������       �      л             �?R       U                 �i3�?~�����>+            �E@S       T                 @��?^n��&�>             9@������������������������       ��mO�H��>             7@������������������������       ��,��H�>              @V       W                  ��?�8+%�#�>             2@������������������������       �                     �?������������������������       �䣣�:��>             1@Y       h                  ��?��G�>�             g@Z       a                 P���?1�XԪ��>~            �_@[       ^                 ���?f�i��g�>t             ]@\       ]                 �p�?@����>r            �\@������������������������       �6chm�y�>F            �Q@������������������������       ��P�>,             F@_       `                 `�X�?C� � �>              @������������������������       �                     �?������������������������       �      ��             �?b       e                 ��;�?�n<�d�>
             $@c       d                 P��?��!t��>             @������������������������       �                     �?������������������������       ���*'��>              @f       g                 ��N�?�.I@�ڒ>             @������������������������       �P�!-91>             @������������������������       ���nӌ>             @i       p                 ��N�?�}m��I�>;            �M@j       m                  ��a?~G9NQ�>
             $@k       l                 ����? ���6��>             @������������������������       � G��̓x>              @������������������������       �                     �?n       o                 @9A�?݉@uk@�>             @������������������������       �;�H�j��>             @������������������������       �      ��             �?q       t                 `s5�?�u�hĞ�>1            �H@r       s                  `%+�?�ܙc�Q�>             @������������������������       ����iO�>              @������������������������       ���J�e��>             @u       v                 ����?�֮Y���>+            �E@������������������������       �                     �?������������������������       �f'~�vQ�>*             E@�t�bh�hhK ��h��R�(KKwKK��h �B�  �态�����o0?u}��{��f���@�T3���L?h��\�W�2�K�S[�?��ثc���Q�-Y?_q+ln�?lJ�s��?M.{�1eS��<<��7U�C���r��N�\p����L�d�?�(1F��@?�i��q�b?3�/H)�d?h����\�?����e�?y1i1�Y�?ެQO=�'?�?�s�f`?�;�l�?��ީ�?���Ō���%�h�;֮>+��?xR�>��D?�9?r�?��-��[?�@Ώ�8?���-W忩DsY�?�\
<m?��] l�?����e�?v���"Z#��9t~i���޸c�UeW�m�<4e���?�Lڮ�?gX��S6ݿ��8�S?�#�1[?�r�I�i?s�oШ_�?�
�`�w�?4����C?@�k�[ݿ��H�b�?�p�"�]�we�?�]�j�?��R-�W忲�n[�/��ճ�*���ۍ�B�3�u�B4?P�|h��P���pɐh������߿��Sׄ������08�pk��P^�|;.A?��?�:��&�T?�!�5�a?e1��o�?�� ;��?������E�Ħ�f_�?�S�C`� �cv �P���$?��+�<��@��E�Gg��?��?��ֿ싀5c��?`Tb8NZ�o���K�e���fYh���tQڍ忼��3�%&�ᒇr�?�[�2��ʿ�]��`�>�i�5�)���u�3l��j�忻'�ʩ���ʿ�uҕL�?�y�8o?uHhtz�?��kwZ�?W~џB�R�Y@U��@f�� k�R'R.a�	c�բ?��t�� V�T�+��[�ʏ<S?�>?@s5�epe?�M6(t~?a�Ps�?�j��?����B?���U�տ��>��p�?^ $���>���i[�[.�j���2�\�Ct_n�1?3!��~z�?�����.�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KEh�hhK ��h��R�(KKE��h��B                          �6Sz?�_�k���>�           �}@                        �lw?Ω�G:g�>           �w@                        �ݤv?~u�R�>z           �w@                        0���?��@���>y           �w@                        �{��?G��W��>v           `w@                        ��>�?��q��>�            �k@������������������������       ����qل�>�             f@������������������������       ��G�>,             F@	       
                 �0;B?���R�>�            @c@������������������������       �q�fs�>o            �[@������������������������       ���̥[U�>+            �E@                        @���?�v�0���>             @                        �V��? �1.3^h>              @������������������������       �                     �?������������������������       �                     �?������������������������       �      ��             �?������������������������       �     ��             �?                        ��6�?�N=I��>             @                        �Q��?�L���>             @                        �/��?@� ��>             @                        �ny?��8��T>              @������������������������       �                     �?������������������������       �      p;             �?������������������������       �                     �?������������������������       �      ��             �?������������������������       �                     �?       (                 ����?�Ҧ�0�>Y            @V@       %                  ��?+��xd�>              @                        8TK�?ڔ�����>             @������������������������       �                     �?       "                 p�,�?�c��Ow>             @        !                 ��~?P����i>             @������������������������       ��Ǎ��)P>              @������������������������       �                     �?#       $                  )5�? *ӭo` >              @������������������������       �                     �?������������������������       �                     �?&       '                 $у�?�&�ύ��>              @������������������������       �                     �?������������������������       �      �;             �?)       8                 �b��?Jy/ے�>Q            @T@*       1                 �� �?#��;���>             =@+       .                 ��;�?�F�'J^�>             9@,       -                 �U�?԰g�ˆ>             7@������������������������       �D���K|>             5@������������������������       ��ϯ�<�n>              @/       0                 
b��?p�%���>              @������������������������       �                     �?������������������������       �      X;             �?2       5                 � �?��c����>             @3       4                  `s�? p��19>              @������������������������       �                     �?������������������������       �      ��             �?6       7                 �p�? jШ]�m>              @������������������������       �                     �?������������������������       �      `�             �?9       >                 ��?��D�RD�>4             J@:       ;                  �_�?��
+;]�>             @������������������������       �                     �?<       =                 H�D�? ��Y�>              @������������������������       �                     �?������������������������       �      0;             �??       B                 �qҍ?oj �<L�>1            �H@@       A                  �?����>             @������������������������       ���7��D>             @������������������������       �      ��             �?C       D                 ���?VWZ_	�>,             F@������������������������       ��|�֮��>             8@������������������������       � ����:�>             4@�t�bh�hhK ��h��R�(KKEKK��h �B(  ����>r������{@
�7;�K�7���|����J�K�?��)&A������I�?N]�6Բ/�9h�ӽ��E��ܿX�N)�B`?���\c�i?c�]��g�?��sFFe�?��T��V�B�sm�?[��(_�d�<�$}vtH�}SB��X�,N'1V�P�	1�4�[��U^/Z忨�i/�b�l���]�?������<��sP^9? �
}��T?��n_�L?<��zL`�?��)O�@E? �px�K?t徏UY�?����p[�? "�7?��5`W�?F`)#W�? �g�?d?۾	-\�?�h�Z�i�?�o�c�3?~{��%mE?�jGj@?8Q���5C?hr+7<Y�?ME�f]�?҂�I�s?�5f)��\�����W�?��:�_Z?����a?��(v�`�?I]5��a�? ��qQ?tX�K\�?ڦ�H�Y�?ޒ�
�?g�P��V��	���o� �3��4?�s�&W�?�
��V�?���X�d)?�}���2H�1�ЀW�?ξ|I�q�#B0���3?GZ�?;WSfG�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K+h�hhK ��h��R�(KK+��h��Bh	         *                  @���?}�$�@·>�           �}@                        �Q]C?��,�EE�>�           p}@                        �0;B?���\��>           Pq@                          �G�?�ݗ\��>           0q@                        �С?��u���>%            �B@                        ��^?c��bB�>             ?@������������������������       �؏*�K��>             @������������������������       �W���>             8@	       
                 0���? �^�12�>             @������������������������       ���}Y�>             @������������������������       �     |�;             �?                        P�}A?�<���I�>�            �m@                        �,$i?B��b'Ҽ>�            @m@������������������������       ��%�ľŹ>�            �b@������������������������       �0����B�>S            �T@                         ��?,`��_�>             @������������������������       ���ca1�>             @������������������������       �                     �?                        0�C�?�Z���>              @������������������������       �                     �?������������������������       �                     �?                        ��,P?�䱲��>�            @h@                        ���I?�k���0�>             ,@                        �B�|?S�=���>             *@                        PX�[?���[�>             &@������������������������       �                     �?������������������������       � Y��S�>
             $@                        .,��?�|��@�>              @������������������������       �                     �?������������������������       �     �i;             �?������������������������       �                     �?        #                 ��� ?u�9���>�            �f@!       "                 xQ�X?�C;LDd>              @������������������������       �                     �?������������������������       �      ��             �?$       '                 ��}?����t��>�            @f@%       &                 �@�?��*�o;�>             5@������������������������       �����@~>             @������������������������       �4F��kI�>             ,@(       )                 gM?伦9��>�            �c@������������������������       ���!<���>             3@������������������������       ���GȊ�>�            @a@������������������������       �     �<             �?�t�bh�hhK ��h��R�(KK+KK��h �BX  ���
�>�d-O�� j<!��?P����}?�x�ơM:�Y\z`2�&�M�=AǬ�縌& �?\�u���Y��T�`�=�U������ ?]�<H�m$?"��}?`��l�?�}KW���^�Z��3�t�e忀7�[*<r?B~��[�?g����?s;4� ����K�E��RL�?��m�H�wG��s��V�?�.߿Z�̀OۭI?��*�]�? �]cfU��c7�Ce忊-t¨��|K���U��+Ԫ�[��M�b�]忠�%CkB�fv��6�8?��`ZY��KJ��?�Pd&Z�!�K�z��9޿������п�����j�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KIh�hhK ��h��R�(KKI��h��B�         (                  �~��?C���w�>�           �}@                        �Zz�?}�Ȭ��>�            �g@                        �S��?O�PQ��>�            �e@                        ��&�?�J��ĸ>�            �e@                        ����?8���e��>�            �b@                        �,�?md��]b�>�            �b@������������������������       �/��3���>s            �\@������������������������       �[
�ҙݦ>!            �@@	       
                 8+	�?PVn\A�>              @������������������������       �                     �?������������������������       �      p;             �?                         <Fm?�� U�>             6@                        @��?��E6�>             1@������������������������       �8�(��ۢ>             0@������������������������       �      �;             �?                        P��?�hA�8r>             @������������������������       �                     �?������������������������       ��S��)�S>             @������������������������       �     ��;             �?                       ��h=�?���Y��>             .@                         @��?ө����>              @������������������������       �                     �?                         �9��?Ҥ�7̀q>             @                         �#�?�-��?>             @������������������������       � @�e ��=              @������������������������       �                     �?                         �g<�?�T�1c�d>             @������������������������       �(j���>              @������������������������       � �)a���=              @       #                 @Q�?#X8.���>             @       "                 P_R�?�W6W�M�>             @        !                  @V��? י�ˏ\>              @������������������������       �                     �?������������������������       �      `�             �?������������������������       �     ��             �?$       '                 �ɡ?p�R5�
C>             @%       &                  �.�?p���,6,>             @������������������������       �                     �?������������������������       ���@�>              @������������������������       �                     �?)       <                 �^��?$~J
�>           �q@*       3                  z�?�F\p�>�            �o@+       2                 ��c�?�!��-�>�            `n@,       /                 ��H�?��W6��>�            @n@-       .                 mu�?�9�o��>�            �l@������������������������       �o��)r��>d             Y@������������������������       �������>�            ``@0       1                 0�Ь?;�;�I�>             &@������������������������       ��elK���>              @������������������������       �*����>	             "@������������������������       �       <             �?4       ;                 p��?����>             (@5       8                 pN�?�����>             &@6       7                 `CE�?@|^�z��>             @������������������������       �P�/-i>              @������������������������       �                     �?9       :                 �j�?���c��>              @������������������������       �                     �?������������������������       ��ۏa�W�>             @������������������������       �      ��             �?=       >                 @���?1K���>             =@������������������������       �                     �??       D                 `V��?��c\�-�>             <@@       A                  ��d�?	�\(�>	             "@������������������������       �                     �?B       C                 0Ɏ�?��~�{�>              @������������������������       ��F���>             @������������������������       ���k�4�>             @E       H                 �h�?+/M�z>             3@F       G                 �j��?c�=��a>             2@������������������������       ���hqj�d>             @������������������������       ��u�o^�<>             (@������������������������       �      �;             �?�t�bh�hhK ��h��R�(KKIKK��h �BH  ^a�b·�@>��#?�Qr��(?t���&?�E�P�X?��^��[?Бq"+�?3�b߀aѿ q?��X?�8��a`�?)��ѪZ�?&R�zFJG?"�;y�N?�8���?'��;f�?��cF����}W�?�H��V���\5�h�?rԵ66�&&�1�AF�ɝ�`�cFBtp?��2D�� G��ǄY���g�X����֮3�iL��V��mX����h.
?�L��	=? �'a>F?�y��&X�?&��i�Y�?�0�4}U忴l��0�Ea%%�
*�|���V�/Q9ѣV����mW忈@�����G����"���8i�F�Ϳ{lJ���:,�$"�zY��S�?��)��xǿ�-�'�j=?L��h�?E66��ӿ·��d�?Ϲ	��Q��^wF}G�I�X�>Y��C���Z�p�,Dd���q8��:�+G���[�?����[��n�_~n忇E�m��3?��9wt�?z��f�?�:mO?�BF��u�?t�i�[6?���,L�?x	#�Z�c����2��h�韸,��n�sX� �TV�zøE�]忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K9h�hhK ��h��R�(KK9��h��Bx         8                  @���?���ݬP�>�           �}@       !                   p��?�@��>�           p}@                        �|_�?��B�>�           �z@                        ЉW�?�bs�
�>�           �x@                        `r�t?lNe:_��>�           x@                        � �J?����k��>E           Pt@������������������������       ����i�g�>           �p@������������������������       ����>8             L@	       
                  9ר?�W���\�><             N@������������������������       �ƌo���>             ?@������������������������       �(p�LQ{>             =@                        ��ݻ?�KI�~�>              @                        �2j?�	�E/�>              @������������������������       �                     �?������������������������       �      Ȼ             �?                        ���?6#�)��>             @������������������������       ������j>              @������������������������       �D�3LhY�>             @                        ��ӹ?9�x�V�>#            �A@                        pM��?� ���>	             "@                         �E�?�P�~��>             @������������������������       ���h�W�F>             @������������������������       �                     �?                        (��?�����=             @������������������������       �                     �?������������������������       � ����w�=             @                        ��4�?<��g���>             :@                        `8�?�3�����>             (@������������������������       � ���jj�>             @������������������������       �^�ݖJ�p>             @                         hTF�?La�I�)`>             ,@������������������������       �                     �?������������������������       �P� �PwM>             *@"       +                 P�bf?�����>+            �E@#       *                 ���?���Z_�>             7@$       '                 ����?��n�ۘ�>             6@%       &                 �t�? ��H��>
             $@������������������������       �{r���t>             @������������������������       ��﬌�S�>             @(       )                 `5�?.(��H>             (@������������������������       � ���%�!>             @������������������������       � ����4>	             "@������������������������       �      �;             �?,       1                 `�Q�?��.t<�>             4@-       0                 ��}?�,>tm�>             @.       /                 ��͎?�M����>              @������������������������       �                     �?������������������������       �      p�             �?������������������������       �      ��             �?2       5                  ���?^�5��>             1@3       4                 ��L�?9O*�_>             @������������������������       ����v�&>              @������������������������       ��r�'1>             @6       7                 f�`?�<e����>             &@������������������������       �8󱽄�>             @������������������������       �
�=a��>             @������������������������       �     %�             �?�t�bh�hhK ��h��R�(KK9KK��h �B�  �\a��$ܾ�A��l��a�<H����"��-���_��mJ �"B�0����\����+�Կ\�@���,?3�y�>�?A}���X�?�X8��[�zD��p�y&~pPf�g��!wo�6�-�qN����Ued�.���<$���%E'4?�k��$�N�>�?�T�v�V��t�jb\�3S�v�O?�B�V�?J��U�?�K����>?(�eN�3I?����T]�?u�1����?��2\j�+?��q�Y�?����V�?��Xe�5?C���?㾀��@��b��9�����U����\快����!?����W�?0��c�U�?�X4��`�?�3$�G?�@<�m�`? $�̿�X?�D��_�?n#'[�?�A��f�?xK�2�??#H��
(�>|���V応��9V�?�Gd�xWH?�;^�?(��ƼZ�?ԫW^jd忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K9h�hhK ��h��R�(KK9��h��Bx         "                 �\/?V�ä�>�           �}@       !                 �}?"O�
�>z            �^@                        �U����c�q�)�>y            @^@                        pF�T?/}����>/            �G@                        ��`?��J-��>             4@                        P��[?�܌�>             (@������������������������       �Ѣ��>             &@������������������������       �      ��             �?	       
                  1�>��T�QG�>              @������������������������       �                     �?������������������������       ���$MF�>             @                        �j��?o���k�>             ;@                        p��v?���}ڰ>             0@������������������������       �#����>             ,@������������������������       �ww����>              @                        ����? �ȶ$��>             &@������������������������       �0�Kگ�>             @������������������������       �`�=���>              @                          ��?c2'��*�>J            �R@                        0~�:?��+��d�>)            �D@                         y��?�5�Ӥ>             ?@������������������������       �!8�u���>             2@������������������������       ���Zn��>             *@                        �p�C?��Aqj�>
             $@������������������������       �\Q�֯��>              @������������������������       ��G@ԙd�>              @                        �-�?:JKFj��>!            �@@                        @B�<?&��3y�>             @������������������������       ��.���`>             @������������������������       ��V��XM>             @                          0�9�?�	�� �>             :@������������������������       �,��Z���>             7@������������������������       � �z瓞�=             @������������������������       �      �;             �?#       *                 P�Y�?��o<s�>^           �u@$       )                 �ڔ�?�\@>��>             @%       &                 �'6;?��I�>	�>             @������������������������       �                     �?'       (                 L��?����h>              @������������������������       �                     �?������������������������       �      �;             �?������������������������       �                     �?+       ,                 �f1�?�iƯ���>Z           �u@������������������������       �                     �?-       2                 ��g?��6���>Y           �u@.       /                 �$I�?q����>             1@������������������������       �                     �?0       1                 ���`?V��x��>             0@������������������������       ��1�/2�>
             $@������������������������       �x�Ӻ&%�>             @3       6                 0��s?ٙ�nѨ>H           �t@4       5                 0Rkz?�{�l�>"             A@������������������������       ���G(^�>             3@������������������������       �Fن�v�>             .@7       8                 �D������N<�>&           `r@������������������������       ��z]�ΰ>o            �[@������������������������       ����A���>�            �f@�t�bh�hhK ��h��R�(KK9KK��h �B�  E�<x��>���Be$?۵���?���ۄ"����� �C�_pI	O�	����S�ؿ�&���j�?i�fY�HW���? Z�?�	5��_��e�^��)?�Jǫ��J?;5��Lp�?�����ֿ��%���F���1Jb忑�aa��ÿ_ |��1?��;��	?WSd�0 �(y?�4�?w�Ĥ�ܿց?ri�D?l[+��տ
���?P���qA?BQm��_�� �c�wW�?lm���W�;����\F?v�Y�Z�?�D��%V�?xl(��s�?^.�:����:�{�QV����ė�L��JǻV��4����T�X#�7\]忏��� [�jQ�D�d�9ϑ���9.��e�?@p#`����X���7?�����h�?�q���%?���>�ڿA�%�*�?�4�3��g�G��:�zڜ�#j�8�?u~�L���딘���?�>ө&�ɿ�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KSh�hhK ��h��R�(KKS��h��B(         2                 �rq?���F	��>�           �}@                        �C
T?�M~���>�            �`@                        �U����ѝ����>U            @U@                         e	a?�=nD�>#            �A@                        P��[?.�
��>             .@                        `��> u|���>             *@������������������������       �                     �?������������������������       ��ו�m��>             (@	       
                 p��3? (�Hg>              @������������������������       �                     �?������������������������       �      ��             �?                         �Sr?<v��ͻ>             4@                        �,$�?2(���3�>             *@������������������������       � �/,0=�>             (@������������������������       �                     �?                        U��?x�L��>             @������������������������       ���竀�>             @������������������������       � �	ļ>              @                         ����?ƞH�3��>2             I@                        �C>?G[#�E�>             9@                        ?Z?^�AGɁ>             ,@������������������������       �                     �?������������������������       �pn4 I@k>             *@                          �P�?&�T�>             &@������������������������       �8���:�>	             "@������������������������       �H��v���>              @                        ���?/��,���>             9@                        ����?"KnU�h�>             8@������������������������       ��h~,�>             6@������������������������       ��M�0�>              @������������������������       �      �;             �?        )                 ����?�:O�?��>0             H@!       (                 `޳?�&欳>*             E@"       %                 8'�?&�V����>)            �D@#       $                 `�ռ?��cH�>'            �C@������������������������       �K�yJ�>             :@������������������������       �̼�yY3�>             *@&       '                 �L+�?�<��P��>              @������������������������       �                     �?������������������������       �      ��             �?������������������������       �      �;             �?*       -                   E(�?p��ZYƂ>             @+       ,                 �K��?h���\Bg>              @������������������������       �                     �?������������������������       �      P�             �?.       1                 Z��?0M��}>             @/       0                 X��?���K��=             @������������������������       �                     �?������������������������       �  ���Sm=              @������������������������       �      �             �?3       B                 `�ہ?&�#cf��>S           0u@4       =                 �9a�?|�s៥�>+            �E@5       <                  ��g�?@����>(             D@6       9                 �u�p?�ۈ�.)�>'            �C@7       8                 l��I?4%%��@�>             @������������������������       �� ��:�>             @������������������������       �N��1�*Y>             @:       ;                   �P�?c��ŉ�>              @@������������������������       �YCڏb�>             2@������������������������       �B'?�u��>             ,@������������������������       �      �;             �?>       A                 �	��? êR���>             @?       @                  �_�?��M�5��>              @������������������������       �                     �?������������������������       �      �;             �?������������������������       �                     �?C       D                 @�q�?w'�8�Ѷ>(           �r@������������������������       �                     �?E       L                 �v��?UQ�>��>'           pr@F       I                 �n0�?HH@yt�>4             J@G       H                 p'v�?(�\J���>/            �G@������������������������       ��'�	��>             &@������������������������       ��q[2�ȼ>$             B@J       K                  ��d�?r����#�>             @������������������������       ��X,�me>             @������������������������       �p����/�>              @M       P                 `�݇?qzd�;�>�            `n@N       O                 �F��?�|����>	             "@������������������������       ����T7��>              @������������������������       �      ��             �?Q       R                 ���`?RǪT2��>�            @m@������������������������       �П�Zg�>              @������������������������       �$�0}X�>�             m@�t�bh�hhK ��h��R�(KKSKK��h �B�  ���#��>�rj}#�ľRUj?�@n0�T??��&n4!�!d���H:?�at�Y忸�*[�3�?g�9�km�H�y�g忙�
�(j�+��Q �N?��wTY?���x`�?�	,m�]忸n���b%����[忓J<9Z�?�k:�-��h*�R%?�Lʵ��.�����Y�??���W忖ǀz�X@?�~x���?	>]*]�?��b�5�A�d�k_L�>�V��f��χv*�?�{��2b�{@���@�-P�D���@f�A�Wꄔ�A>�e���|ȿ���&]�~�� a�yv��Y�Vh�c�g�It�th���:$? Tk eE?,;
Z�?�ju�W�?�/�S��-������d�VY�U���SV�8Y�~zU��<�R�?Jaɏg�>?.�]m�\2?!v����*?�M/���O?|��N^�?72�.W�?�o�Qi&?|8���?��PG��տ�dzNg�?U����h? G'�l?��\�jf�?E�e�j�?�ˉ=_�? ���c��>��/�k忤7!����>A����2�����i%�I)���ڿH�Ɏ�?����U�dx�u�Z��(H�@b�y���$I?�j�gQ?�G� �?aE�Wun�?��Y~�?�-+)`�?�΁���?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KCh�hhK ��h��R�(KKC��h��B�                           P��?�$y�u�>�           �}@                        ����?�lzF4�>�            `f@                        �r�?�Rtn��>�            �e@                        йϷ?=�ᐒ>W            �U@                        ��6�?k:�o��>Q            @T@                        0gç?!@�^�-Z>N            �S@������������������������       �,kN��'>G            �Q@������������������������       ��#)���>             @	       
                 �*c?5
Y8��>             @������������������������       � .	-�>              @������������������������       �      �;             �?                        ���?0����>             @                        0���?����B�>             @������������������������       ������>             @������������������������       � ��6�MQ>              @������������������������       �                     �?                        p�Ӄ?�vM���>X             V@������������������������       �                     �?                         ���/�����>W            �U@                        ��/�?��-!]@�>             9@������������������������       �/�rZ���>             *@������������������������       ����#u��>             (@                        �Q�?�Т�Y�>>             O@������������������������       �                     �?������������������������       �fDjT�>=            �N@                         `���?�)���>             @                        0�!�?@���E�>              @������������������������       �                     �?������������������������       �      �;             �?                        �Ч?�����j>              @������������������������       �                     �?������������������������       �     �7�             �?!       &                 ��?S9.��>%           Pr@"       #                 X椐?������>             @������������������������       �                     �?$       %                 �w�?;a�9*��>              @������������������������       �                     �?������������������������       �      :;             �?'       4                 p��?�2@�¡>"            r@(       /                 `]P�?�"d��>�            @n@)       ,                 ;�?�d�VhQ�>�            �g@*       +                 �&��?�ҿ��9�>|             _@������������������������       �â3��O�>z            �^@������������������������       �Sh��m��>              @-       .                  ^M�?텑��a�>B            �P@������������������������       ��̧���>#            �A@������������������������       ���M=*��>             ?@0       1                 ���?]�͆4�>4             J@������������������������       �                     �?2       3                 �y��?d`��!A�>3            �I@������������������������       ��0X��.�>/            �G@������������������������       �����>             @5       <                  ��?��sŮ@�>0             H@6       9                  ��?#F��$��>             @7       8                 ���?!L^�>             @������������������������       �                     �?������������������������       ����3��z>             @:       ;                 ����?6�8~��T>             @������������������������       �fd�}Y >              @������������������������       �                     �?=       @                 pg��?����1x>)            �D@>       ?                 �'��?�C>��5>              @������������������������       �                     �?������������������������       �      P;             �?A       B                 xE�s?Ė(��t>'            �C@������������������������       ��\�|(Q>             4@������������������������       �<�آz>             3@�t�bh�hhK ��h��R�(KKCKK��h �B  .�-B�Ǿ�;j��?��k�C�?�i�$V����`Y��e�0g�G:��^|�	����\�r�6ʑS?H�H�V�,�!�Zk�?��`�mFE�A���6�x���U�>�iP�Y�nWF�Aa�����T�0?�F��e�?�BQL�-?��$�	7D?j �����U=FTF��?�)u���?9e,]��!�i�?���`f�N�\�����a��˱d�L]��4^� @3a{�1?Dk��	X�?��]ȗU�?;%�X1	�E����sR���[�/l� о�_�9?���Z�Y�?\=��tU�?C(c`X�3����%�P�+�r�!�J�ߌ
�=U4�̿U�M��o�?~p*?��3��jYY�⿚���r㢿
?��bS ?{����e�?crK�?��3�`��?wIKt�h>ݩ(?֗�t.R? �\��_?	�b�&W�?�L�c�?51
��羱ʒ	�U�?����oV���{u��>��R9��A�q��M�W�fn�ðX�՗�4�b?�џ+�V�?��U��̿�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K]h�hhK ��h��R�(KK]��h��BX         6                  �=�?�7U4Q�>�           �}@                        ��{�?s)�[4
�>            q@                        ��p�?̦�O@��>�            �m@                        ��'j?�y�	�f�>�            @l@                        �<�?Pχ/\�>�            `d@                        pb!i?_�2�ԕ>�             b@������������������������       �s�tȏ�>[            �V@������������������������       �Qb�U�>6             K@	       
                 0Ԃ�?�u�a��>             2@������������������������       ����#��>             *@������������������������       �Z�N�>             @                        `�Q�?�&�Zݢ>?            �O@                        �p�?�P��L�>+            �E@������������������������       �]�ێ��>             7@������������������������       ��[.�&�>             4@                        �+�?>d��>             4@������������������������       �h�DZ�>
             $@������������������������       �7@��>
             $@                         P���?����a��>             (@                        ��Y�?]���cp�>	             "@                        8��?�/��q>             @������������������������       ��(Fo+>              @������������������������       �                     �?                         ���?0��\k�}>             @������������������������       ��8wC4u>             @������������������������       � B=��6>              @                         ��?s�{�K�>             @                        P$��?T��+I�>              @������������������������       �                     �?������������������������       �       �             �?������������������������       �                     �?        '                 0vb�?�6�X�>$             B@!       "                  ��~�?�%Z��>             *@������������������������       �                     �?#       $                 �͡�?���!�]>             (@������������������������       �                     �?%       &                   ���?����N>             &@������������������������       ���'�A�Q>             @������������������������       �^�I�7,>             @(       /                 `횃?�,V%�e�>             7@)       ,                 p��=?>`y�E��>              @*       +                 @��?�f{��>             @������������������������       �                     �?������������������������       � iKp�=             @-       .                   ���?�|���l>             @������������������������       � ���,h>              @������������������������       � ��
�I>              @0       3                  0p��?�ڗ���>             .@1       2                 tم�?|䌼��u>             *@������������������������       �*(_�n>             (@������������������������       �                     �?4       5                    �?``���n>              @������������������������       �                     �?������������������������       �                     �?7       L                 `7S�?��'�.��>�            �h@8       E                 ����?���'�V�>             0@9       @                 �ڡ3?�Q����>             (@:       =                 ��jm?���}}>             @;       <                  �j?��?_e>             @������������������������       �@Ob5�|N>              @������������������������       �      t;             �?>       ?                 ��q~?PR
��6W>              @������������������������       �                     �?������������������������       �      ;             �?A       B                 �ڡC?*���
s>             @������������������������       �                     �?C       D                  `S��?WaL�G1>             @������������������������       �                     �?������������������������       �j�t'�*>             @F       K                  ����?r�@�>             @G       H                 @ϡ?��{>�>             @������������������������       �                     �?I       J                 �Zv�?�"]��Hq>              @������������������������       �                     �?������������������������       �                     �?������������������������       �      ��             �?M       P                 @�Dv?�He��<�>�            �f@N       O                 ���@?���39ɵ>              @������������������������       �                     �?������������������������       �     �z;             �?Q       V                 ��/�?�=��Y��>�            �f@R       U                  ���?T81@��>             @S       T                  P���?��.]�_^>             @������������������������       � ���<>              @������������������������       �      `�             �?������������������������       �      M;             �?W       Z                 �p��?6����Ζ>�             f@X       Y                 �W�?f��P^x�>             @������������������������       ������l>             @������������������������       �����dk>              @[       \                 `�ޮ?-�&�>�             e@������������������������       �������>             @������������������������       ������>�            �d@�t�bh�hhK ��h��R�(KK]KK��h �B�  �+#t��>6'k���?�ۻe�>S&���?�������u���?�� ��:+�?��{�?�ֿ�8���6?Й�.�O�?Jg����?�+*)0?z�c�(?a0 �:��?�y��g�ɿ��/��B?���ϑ�?W�3A�$�?�~��UtA��5zNcJ�xœ�@j+?��Q����?��cX�?����U��T�9�[���\^忘T��(�2?�:۫f�)U��YU��`���U�ѱ[�_Z�?�x��9?��"M8��<'6o�[�?�ռPv&�L�VqX���v�5V!��T��V忊m�f�U��� [~E? �v=-�U? �)JtG?S�H�;^�?;��W�?�PXs5p_?��Ya�?��<��^�?it��3?e��pd)?^u��%�?��iE~W� �C�;�P?��/\�?1���Y�?�T(�h���o��=��f
�)�+��14�*@B�8�`65�I��֔�_Z�0�IX���ŕlB,�ܴ�PW忆[3�U忡QV7� ?�2�F�X�?�UF�io�����iV��o꫻U�z��O\S��+���F��4,xU�+���ROP��/*\忐�$cY�_�J�-d�˄��S���ȑ0*WR?M&���a�?��6xqU�T^�J�K�v�|.ʰF?U!��l6O?ocW,[�?��p�XY�?\���U忎N����
2468
B��;	��W忞\�v@]�������>�����?F��:�H˿�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kch�hhK ��h��R�(KKc��h��B�         4                 P�$�?��h��>�           �}@       !                 ��{�?��Hu��>�           �y@                        0���?ҖvĀ��>�           Px@                        ��a,?����L�>O           �t@                         �Y�?	QN/�;�>�            �d@                        �&Ұ?B����(�>�            `c@������������������������       �;�����>l             [@������������������������       �lٮm�a�>/            �G@	       
                 ��o�?�_@��>
             $@������������������������       �                     �?������������������������       �;;���%}>	             "@                        0	q?A}UHy�>�            @e@                        �rq?,i���T�>j            �Z@������������������������       �w�9�*��>+            �E@������������������������       ����uw�>?            �O@                         p%+�?��1Zkr>@             P@������������������������       �                     �?������������������������       �p��%��o>?            �O@                        ��?��o�욤>6             K@                        .�X?���:�>             ;@                        p?�����R�>             &@������������������������       ��K�Pa�>             @������������������������       � R�rA�V>             @                        P�$�?���}>             0@������������������������       �`�~ʦ�]>             @������������������������       ��MG�FSv>             *@                         ��?��R��>             ;@                         ���?����>             2@������������������������       ��� b�>             &@������������������������       �����>             @                         ࡑ?���+��>	             "@������������������������       �                     �?������������������������       �\�pO�<x>              @"       +                 ��N�?��`��K�>             9@#       *                 ���?a4�9��>             0@$       '                  �t�?!�b�匭>             .@%       &                 �W�?��<�i�>             @������������������������       ��ЍҮ�>             @������������������������       � �v�Vly>             @(       )                 ،��?�s��e��>              @������������������������       ��z�^E��>             @������������������������       ���ɋ���>             @������������������������       �      �;             �?,       -                  ���?�-���ñ>	             "@������������������������       �                     �?.       1                  `���?��_���>              @/       0                  s��?x���Q�>             @������������������������       �@��B�*>              @������������������������       �                     �?2       3                 ��&�?��5&?>             @������������������������       � ���~�=              @������������������������       ���_��>             @5       L                 P���?P~=���>:             M@6       C                 ����?z[O6e�>             =@7       <                 ��c�?�xZs֘>             8@8       9                 ��D?�6��C�>             1@������������������������       �                     �?:       ;                 8蠂?���ӑ��>             0@������������������������       �ܮ{�N҄>             @������������������������       ��ݫ]!Uz>             (@=       @                  Џ~�?J7ֺ�Ӡ>             @>       ?                 �j%?.��}��x>              @������������������������       �                     �?������������������������       �                     �?A       B                 ����?H;J���>             @������������������������       � +b�n>             @������������������������       �     ��;             �?D       G                 (tns?9�#��u>             @E       F                 {��?��@^�;X>              @������������������������       �                     �?������������������������       �      P;             �?H       K                 `'v�?��$�D>             @I       J                  0B�?�3�i�8�=              @������������������������       �                     �?������������������������       �      �:             �?������������������������       �                     �?M       X                   ��?Z<���>             =@N       U                  ����?/Κy�ǐ>             2@O       R                 �@�?�!�~}�x>             0@P       Q                 06y?2�s�ij>             ,@������������������������       �                     �?������������������������       ��	Wa��b>             *@S       T                 ����?p���
�d>              @������������������������       �                     �?������������������������       �      @�             �?V       W                    �?��Y�{��>              @������������������������       �                     �?������������������������       �      `;             �?Y       ^                 ��f?�A@��4�>             &@Z       [                 0I��?P�����>             @������������������������       �                     �?\       ]                 ���H?�ꜧ��a>              @������������������������       �                     �?������������������������       �                     �?_       `                  ���?垤�� �>              @������������������������       �                     �?a       b                 �C�?ڞku��=>             @������������������������       ���M�o�=             @������������������������       � ���#>             @�t�bh�hhK ��h��R�(KKcKK��h �B  c�n׾I5u��>V��������4�>Ջ{p'��8�I�{�����~���A�g�ϿfZ���<:?��Y�g�?O$*_m��?̴2�1S?�:^�a\'?R���.��*lkOI��?Pr��e��2�)Z��A3�տSc%ڙ�*���ע�B�!�ǽ��N��D1��#ٿ����._��z��:$4��ÎKvY��9U��X�m�Q�Wy$?�[�U�:?����A�?�Qz�`���ZJ,47���@\忬30?�X忤Y ;aE?�!_��}Q?t�H
�3L?�w���aW?���Ӣa�?��G<!Y�?s�k��7?� '�/̿Sǈt
[�?��Ѣ5l�?ˠ��r�t��	ob�ef�ؔ*? ����G?(-Q|*V�?����_�?�դ�����}�V�=ս�U���V���'�h��K�;���x���A�^�fS��6�1��ݏW�?�Q2e�9���ɏZ�ؚ����z���v�P����pY7��`֞U忷����X�B�w$NEU��kB I^��X�3�U�j��t0&? x��5@?6?�7W�?�����X�?��!�����>���w��dL�c�U�.1gU応�DF�U���T/e?֒%� "���qHD˾�P/�&?���TX�?��tW�8�?l�k�{B�����|Y�L�rXW��h#]��S����z^�ٙ�_lY�0Ne'�9? ��w��R?~pS�^�? �J�:L?G�PY�?S-�1[�?�!m�?,9��]�?(9�����?lU��O��MV忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KWh�hhK ��h��R�(KKW��h��B         8                   Y��?f>P;���>�           �}@                        ��0b?�,�Б>�           �y@                        0�B�?fX|X~
�>�            �i@       	                 �K��?k_MLC%�>�            �f@                        ��+a?Ҕk=̓>�            `f@                        p'v�?U�+���>�            @f@������������������������       �B[I�:`�>i            @Z@������������������������       �|(b6!�>I            @R@������������������������       �     �λ             �?
                         �a�?���M��>              @������������������������       �                     �?������������������������       �                     �?                        �6�?��f2ff�>             8@                        P���?J(�2m��>             @                        ��0�?a���~�>             @������������������������       ��K����c>              @������������������������       �����BGv>             @������������������������       �                     �?                         �9��?�YC1i��>             1@                        8�#�?ԅ�lɦr>             @������������������������       � 9�GO>             @������������������������       �      4�             �?                        �~+�?�o,@�>             *@������������������������       �                     �?������������������������       �F��$.?i>             (@       )                 �D���(ʍR�>�             j@       "                   s��?i�[�^�>I            @R@                         P��?"H�&�[>             ?@                         ��?��Hwr�)>             :@������������������������       ������>              @������������������������       �
D��ϣ>             8@        !                 �,^�?��&�K�|>             @������������������������       �                     �?������������������������       �|��l��D>             @#       &                 �1��?'e�yQ��>*             E@$       %                 @K<�?�fl;3߄>!            �@@������������������������       �*�N��tZ>             9@������������������������       �	�pCM�>              @'       (                 ����?�C$�>	             "@������������������������       ���X��Ip>             @������������������������       ��[�F>�\>             @*       1                  �g<�?Ց�TU��>�             a@+       .                 n~?�f@�s>+            �E@,       -                 p�n�?7��Zs>              @@������������������������       �����X�a>             7@������������������������       �J��3(u>	             "@/       0                 ����?Џv/0>             &@������������������������       ��$��w>             @������������������������       �Q�Xw�n&>             @2       5                 0%�9?�T'� :�>]            @W@3       4                 ��0�?����>             @������������������������       � ��ɫ�L>             @������������������������       ��evKl�>             @6       7                  ���?�!�Z�l�>V            �U@������������������������       �L�By�(�>3            �I@������������������������       �T ���!�>#            �A@9       B                 0�Z|?��� >�>:             M@:       A                 �vq?A@��L+�>             @;       @                 PT�\?����wb>             @<       =                  0�9�?������=             @������������������������       �                     �?>       ?                 ��ue?�OI�e�=             @������������������������       �@Ҙ��K=              @������������������������       �      ��             �?������������������������       �      @;             �?������������������������       �                     �?C       R                 �2*�?n���>4             J@D       K                 T�Y?׃�G��>1            �H@E       H                   p��?DO��+Ѓ>             8@F       G                 p�l�?�m1��>             @������������������������       ��t.k�U>             @������������������������       � �K��Wc>              @I       J                  @���?n��fG�`>             3@������������������������       ��` ���I>             2@������������������������       �                     �?L       O                 `�Q�?���L�Cx>             9@M       N                 (�i<?=��~��>             @������������������������       �                     �?������������������������       � xT�Ⱦ�=              @P       Q                 �=�?��#��h>             6@������������������������       ��V��v>
             $@������������������������       �Q��(}>             (@S       V                  �u��?R"�����>             @T       U                 `'v�?~�\�NQ>              @������������������������       �                     �?������������������������       �      �             �?������������������������       �                     �?�t�bh�hhK ��h��R�(KKWKK��h �B�  x
`�6�>C����Q��H�>ל/w���kcwm���9Z��@��yV�?P
%RY"ܿ<��m$[�?6�^�*�S?G��wU�2�<�b�?�wZԳ6?��C�&�P?>�>\sE?��8f�p���T.[�?�JF�jg�?x_�_7�?I��</AB�h�yAY忰��;V� �i�1?F�PNb]�?�<�0�W�?bp���E���
+�xI`<��N�c�m!��sdcV忙����U�bc$?d���Y�?Ykl>����2��z�a6�/�s(H�-�y�!W��\<�]�܃$O�I�~��C9[��i�X�*�\a��>g�sn;_!��B�r�+��P	�������X�х�>�?���*V�?�+��U�?����6�?��jI?b}Σ�V念��r�c�?�;�m?�ة���?����O_ѿ3�_(��!?t�����G?���5�����3F�r��{U�ٰ4P�xɾ9HS�VU忹;�h_U�� ���W�K('p�?�1��*?}�{"!p�>?�p���#�����B��Bi����E�&�\�A�v ���Gw�;�����z�w�X�G�6*?���JG?�G�a�[�?�\�W�?�V��/!?~�Q�G�?c�5��U�? T�w�E? ��k�u#?9���V�?��EjsU�?Lڤ��^�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K1h�hhK ��h��R�(KK1��h��B�
         0                  @���?�NCG�>�           �}@                         ��^�?j��!�>�           p}@                         ys8?pq�>���>             1@                        `7p.?D2/B��>              @                        �9=h?��*����>             @                           �?h�Л`�n>             @������������������������       �YJ!�X>             @������������������������       � 2i>              @	       
                 (�ȓ?��A��|>              @������������������������       �                     �?������������������������       �      P;             �?������������������������       �                     �?                        �fA?���sZ{>	             "@������������������������       �                     �?                        Ƚ�e?�F�5f>              @������������������������       �                     �?                        ��XD?���jܠM>             @������������������������       �                     �?������������������������       ��?��]b?>             @       #                  �=�?����>�           `|@                        `��?��`��>           @p@                        ��IL?��OV��>�             h@                        ���J?2�TQr�>
             $@������������������������       ���n��>	             "@������������������������       �                     �?                         sR?�=���>�            �f@������������������������       �ĩX�Z�Y>
             $@������������������������       ���Z$��>�            �e@                         Ш��?�X���^�>C            �P@                         @V��?�4��7>              @������������������������       �                     �?������������������������       �                     �?!       "                 p��?"pV��V�>A            @P@������������������������       ��h`��>             6@������������������������       �c� ^f�>+            �E@$       )                  Ɵ�?i50Ú�>�            @h@%       (                  �J�?��h��>P             T@&       '                 �.�x?J6�W{>O            �S@������������������������       �c�����>             @������������������������       ���&(�t>K            �R@������������������������       �      ��             �?*       -                 �B�?��k6��>r            �\@+       ,                  P?��?(i�S��>              @������������������������       �                     �?������������������������       �                     �?.       /                 p���?�f�	��x>p             \@������������������������       �@�r�)L�>             @������������������������       �n1t�ov>j            �Z@������������������������       �     ���             �?�t�bh�hhK ��h��R�(KK1KK��h �B�  O�K��Ӿ�.>��۾������)�eo�Q��A�7˨�1�4�'�vv"��k��
2�?#6)�`W�f7�9�J��F���[��0.��W��Tc�`快�ç�?�*½�Y�?�����Q�>�7���W�?)I��l����bD?V�?���DV�?||C��>���GB?D!O���>�"�TF4?�`�f�1�?zA��]�?��8���N��W���c��u?��Oa�w ? \,I?>���Y�?RѪ�Y�?�1(�x�?��2 ���	��G���? ����D����+���ٛ��x���gژ]������Ϳ�}~1�`忍�!v`�> *�jW?K���X�?��VR�a�?�k��E�� 3�{�����Y������Y�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KIh�hhK ��h��R�(KKI��h��B�                           ��^�?�����>�           �}@                         ys8?�LUsC}�>             1@                        `7p.?CZ|�"��>              @                        �9=h?VҀ�ƅ>             @                           �?�v.%n>             @                        �Ls?s��V>             @������������������������       �                     �?������������������������       ���,�2>              @	       
                 �vQ? ���-��=              @������������������������       �                     �?������������������������       �      @;             �?                        ��?����{>              @������������������������       �                     �?������������������������       �      P�             �?������������������������       �                     �?                        �fA?,���{>	             "@������������������������       �                     �?                        Ƚ�e?�|�zL�d>              @������������������������       �                     �?                        �$I�?P����dQ>             @                       f6?�?t/����?>             @������������������������       �                     �?������������������������       ����џ�3>             @                        8�K�?p#�� 3:>              @������������������������       �                     �?������������������������       �     ��:             �?       8                  ����? ���O�>�           p|@       )                  �_�?����-�>           �p@       "                 �\ͥ?P92wێ>R            �T@                        ��IL?�rF[㕕>             6@������������������������       �                     �?        !                 �2OV?R�f�>             5@������������������������       ���^v�>             2@������������������������       ���Ͽ.�>             @#       &                 ��_�?f* �$u�><             N@$       %                   Mt?#����Q�>:             M@������������������������       �����{>             ;@������������������������       ��/f9��>             ?@'       (               �$���?��ӑc�O>              @������������������������       �                     �?������������������������       �      P;             �?*       1                 �C8�?�$����>�            �g@+       .                 r�4?��J�O�>1            �H@,       -                  .:q?눝�J�>             &@������������������������       ���YǷ�>             @������������������������       �)o�z��`>             @/       0                 P��?��bҕ>&             C@������������������������       ��Q�g�>             =@������������������������       ���G��P>	             "@2       5                 pTF�?�?ӌ>�            `a@3       4                  �j%?@R���z{>             @������������������������       �pb?o{>             @������������������������       �����->              @6       7                   ���?��ܘ��>�            �`@������������������������       �r����>r            �\@������������������������       �,�����>             4@9       H                 ��]�?�vw���>�             g@:       A                 �e�?��&<[�>�             g@;       >                 �I��?�Ȁ�n�>p             \@<       =                 @�N�?������>g            �Y@������������������������       ��9�8j~�>`             X@������������������������       �B	����>             @?       @                 (�t�?�����ʖ>	             "@������������������������       �                     �?������������������������       �_|r�B�>              @B       E                 �Ö�?򾬧�Շ>H             R@C       D                 pO�v?�;.\'B�>	             "@������������������������       ����X��>             @������������������������       ��|��U�>             @F       G                  (��?P\��d{>?            �O@������������������������       ��}u���>!            �@@������������������������       ��PuB�c6>             >@������������������������       �      ��             �?�t�bh�hhK ��h��R�(KKIKK��h �BH  70m���>I��fP-?@�}$	�B?H�Tk�x6?����#?�j.�9��M\�Q>V�?��+V� ��@ �:?�`ҒW�?�m���W�? V�IK?���[�?��CX�?���aa�?\y�����|�~�Y��wx��>�Xވ�W�6�r��9?�yF��!?��$�V�?��� V�?E��\����J=5V�s���ZU�q�����۾�n|����[ȵ3GY?�ئM{�����[]����3 �UMc]�>Կ�3�ES/�?'y�d)8 ?̎��n#?,��"0��?V���H�?���ì�@��#B��X�鸧�qW��W:jI#�(���A.�cQJ(s-?������?��/�KW�s�G�/�7����]z�o�}b�Լ?\�p�9�����lZ*G?m�غZ�?���W�?�ϛ�����>ލC���`�:�f��$����?�f{�?>Jh;(�>\�e'�I?�����
e�}�Y����?��/z�W@�\#���_�AY��r��i
wͮ?��B/��A?L�5}�\�?�6�JGɢ?xR�?bl]>�?H���!V心	��Z忔t�bub�      h,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KMh�hhK ��h��R�(KKM��h��B�         4                 �)�?������z>�           �}@                         ��?-���z>�           �|@                        �rq?e�>��e>�            `j@                        p���?��>��a>�            �`@                        ��gn?^X��dX>�             `@                        ����?�P��M>{            �^@������������������������       �$��mV�F>x             ^@������������������������       ��!v]gWx>             @	       
                    �?7��mI�>             @������������������������       ��2x"FA>             @������������������������       �                     �?                           �?j���I�>             @������������������������       �                     �?                        ��>?�+�h�YZ>             @������������������������       �                     �?������������������������       ��t��_">              @                        0�Q�?��֟��j>O            �S@������������������������       �                     �?                        `s5�?�gu+g>N            �S@                           �?�6@U�{�>              @������������������������       �                     �?������������������������       �     �O�             �?                        p=N�?Q��c�`>L             S@������������������������       ��q+�(]>K            �R@������������������������       �      `�             �?       %                 ��Zy?m���>�             o@       "                  �x?cv�:�P�>             3@                        ��=�?/��ai�b>             1@                          ���?��_��\=>             .@������������������������       �z�2�[�/>             (@������������������������       � {��G�$>             @        !                 ��?�j�t��v>              @������������������������       �                     �?������������������������       �      ,�             �?#       $                  ����? UwsnT>              @������������������������       �                     �?������������������������       �                     �?&       -                 P8��?�%1�mH�>�            �l@'       *                 �r�?&B�ϵ��><             N@(       )                 @=��?�֔j���>              @������������������������       �                     �?������������������������       �      X;             �?+       ,                 �^9�?�g:~b�>:             M@������������������������       ��wQ�<��>             :@������������������������       ��֧Y�^�>              @@.       1                 0I��?��,�q>�             e@/       0                 �ȿ�?�I�M儀>             @������������������������       ���S(�Z>             @������������������������       �      p�             �?2       3                 �6SZ?��[�Zo>�            @d@������������������������       ��xb�r>f            �Y@������������������������       �s�F@a�b><             N@5       :                 p�ռ?ْ��Rw>             *@6       9                 �kS�?��!Ț�k>             @7       8                 `s5�?�Qs;�$P>              @������������������������       �                     �?������������������������       �                     �?������������������������       �      `�             �?;       @                 ����?f�0�)>
             $@<       =                 ��>�?�D��>             @������������������������       �                     �?>       ?                 ����? \�S��=              @������������������������       �                     �?������������������������       �       �             �?A       F                  �x��?3X�i*>             @B       E                 Љ��?�<�B�=             @C       D                  ����?�y�=�=              @������������������������       �                     �?������������������������       �      �             �?������������������������       �      �             �?G       J                 ;��?�]dc���=             @H       I                  ���? �Z�'�=              @������������������������       �                     �?������������������������       �                     �?K       L                  ��^�? 6z
:K�=              @������������������������       �                     �?������������������������       �      �:             �?�t�bh�hhK ��h��R�(KKMKK��h �Bh  ���+���>,�⤯I��1U�:��٘�����>w���/㾊��5���;KY�t�ڿ]�{o��?��� A0?�[	j~��?%�>�([�?j�S\�":?�?��[�?a�܈�#?��X�TW�?������?����A�셢��Y���C���t���5=?*�TZ�?���uuU�.����2��o����vl)X�?4������>����+?^pR�8��,�0n���y����fV� ��V7?�HW��X�?���~�U�? R�$�%a?Ԗװ�a�?��Z`�?�D�B�>]h�G?��0h�<Q?'���:b�?�;7�V忤\���?����`�?;���x�̿(4�Jv(������B�1��w�!/��k�0@[忨%u���g�I�qǿV��i�?�?��zSs�&?U��;�E? ġ�H�@?���6�X�?@��zW�?U@�Z�?ah@=c�>�����^?a\(�vU�?  5��?�`��U�?�X�U�?���V�>A^������/°���n|�"~U忁��ёU�U���U� �o�"?  XE�C�>�
�/rU�?i ŅvU�? �3>Ux?�����U�?iG5�U�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K9h�hhK ��h��R�(KK9��h��Bx         0                  @��?p���cx>�           �}@                        �\/?����:x>�           0}@                        ��S�?r
���z>y            @^@                        �xK�?a���N'y>_            �W@                        �=E?g"q�v>[            �V@                          �G�?1=���w>K            �R@������������������������       ���S�S$p>             1@������������������������       ���sn�w>:             M@	       
                 @�?���_f>             0@������������������������       �GP�j�T>             .@������������������������       �                     �?                         b��>�`���`u>             @                        ��g?����Μ4>             @������������������������       � ���i�=              @������������������������       �      p�             �?������������������������       �      G�             �?                        @�?�#���z>             :@������������������������       �                     �?                        жd|?7��Ev>             9@                         �tx?�}�6�qm>             4@������������������������       ��	�_.d>             3@������������������������       �      p�             �?                        ��`�?"t��]�~>             @������������������������       ���H�[>             @������������������������       �      H;             �?       !                 P�Y�?���2�w>Z           �u@                          ���?:I�q��~>             @                         �.�?0��{zU>             @������������������������       �                     �?                        ��N�?��V���>              @������������������������       �                     �?������������������������       �      0�             �?������������������������       �                     �?"       )                 �/��?ӏK�vv>V           `u@#       &                 ��{�?'��Y��u>*           �r@$       %                 0S�r?�L*#�Ot>
           �p@������������������������       ��Si�y>p             \@������������������������       ��*3?�o>�            @c@'       (                 ��N�?p4_
�#}>              @@������������������������       �y��n���>             4@������������������������       ��Y�5z`a>             (@*       -                 ��F?KG��a�z>,             F@+       ,                 @��8?����ۅ>             6@������������������������       �����,�>             3@������������������������       �$�ļv>             @.       /                 � �J?�`�)�E>             6@������������������������       �                     �?������������������������       ��Z-y�B>             5@1       8                ��#+y?��3]�u>             @2       7                  @���?��Z�3�`>             @3       4                �}��?T���5;$>             @������������������������       �                     �?5       6                  ��u�?�dO���=              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �      `;             �?�t�bh�hhK ��h��R�(KK9KK��h �B�  5�����ݾ;Y�IY���U�u��?Y5C&����S��6�&�>�V�7�	?=�d$�Cֿ�Ԡ5A��?�TT]u �-i�Uڿ��2GY�\ ����<��F�C�%ZhZX�(�v�"Y��%��U�? *�/�B%?�nÅ!Z�?|Ȋ9��!?��~}Rf?�/D�;�?8_�>X�^ \`9?�d�X�?���V忠?��~a��A��M�=�e�TZB"1�J'�U��S�/�7�ɴ�{W�s��aW� �	�Z�O#�C�>��8��;L��*=c�������5ɿ�|D�?�xMvh��i!aܿ��Ep��?.h�psK?)�Yy'?�S��f��?�Y�Y�?��}������{��V�������^��S80?kVrU� ?�;Qa]�>����U�?'e�4�;Ҿ�Ȑ�VU忯��9`U忶g�Y�W�?����FY�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kch�hhK ��h��R�(KKc��h��B�         8                 P�$�?S�����~>�           �}@       !                 ��{�?5���7�>�           �y@                          �G�?-�>�           Px@                        Pz�? Ɇ��r{>3            �I@                        ��H�?�8�j�x>$             B@                        ���s?`�*�
v>"             A@������������������������       ��`��efc>             ,@������������������������       ��q��Rw>             4@	       
                 ���m?0�ZmiE>              @������������������������       �                     �?������������������������       �      P;             �?                        p(�?�s����u>             .@                        �Hw�? ����@>             @������������������������       � ���J>              @������������������������       �                     �?                        �D�A?�"�V=�f>             (@������������������������       ���wh9t>             @������������������������       ���Ɏ�?>              @                         �P��?o
7$Z>R            u@                        � �8?�n�E�z>;            �M@                        0��\?�SW���{>*             E@������������������������       ��t� �)r>             8@������������������������       �8�xl�}>             2@                        ���?j��,l>             1@������������������������       ���D(�a>             .@������������������������       �0�C���j>              @                          \��?���
w�>           pq@                        ��]�?w�f�{��>	             "@������������������������       �ພ�k�h>             @������������������������       �����>              @                            �?���W>           �p@������������������������       ��f|��>�            �b@������������������������       ��Ij*�}>y            @^@"       /                 �Z#�?X��1�>             9@#       *                  �t�?�k��$$z>             4@$       '                 �W�?~��N)St>             @%       &                 `U�? �Y�hVV>             @������������������������       �                     �?������������������������       � �[�^7>              @(       )                 ����?�cكT>             @������������������������       �T�2C�<>              @������������������������       �      0;             �?+       ,                 p\C�?S�i�7r>             ,@������������������������       �                     �?-       .                 @���?��9�o>             *@������������������������       ��nᆂb>             @������������������������       �)���0�k>             @0       7                 `��?�zX���>             @1       4                 A��?Ƣ�t>             @2       3                    �? ;V�%>              @������������������������       �                     �?������������������������       �                     �?5       6                 0���?�$q.\�=              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?9       N                 ��F?�&�5wp>:             M@:       I                 ��q�?zhz��s>             ?@;       B                 �(�?j���V�p>             <@<       ?                 0*��?���(�oR>
             $@=       >                   ��?`cE��U>              @������������������������       �                     �?������������������������       �                     �?@       A                 \��X?3�Ib8>              @������������������������       ��A�<��=              @������������������������       ���i fJ>             @C       F                 �b'�?v��T�Ir>             2@D       E                 p�V�?��ٰ0�o>             (@������������������������       ��6&<�`>             @������������������������       ��P��"�c>              @G       H                 �2*�?Ħ�cc>             @������������������������       �w���V�U>             @������������������������       �p�*��6>              @J       M                 ����?L���[>             @K       L                   u�? �F�YT/>              @������������������������       �                     �?������������������������       �      0�             �?������������������������       �     �;             �?O       V                 ��!�?�py�'`>             ;@P       U                 ��?��+�3zD>             @Q       R                 ��d?�Шr�8>             @������������������������       �                     �?S       T                ���?�r�z�>             @������������������������       �                     �?������������������������       ���q�_��=             @������������������������       �      0;             �?W       \                 �s�?�C���`>             5@X       [                 �I�?�>��+�h>             (@Y       Z                 �מp?�#X�S>             &@������������������������       �
[�2�WR>             @������������������������       �38��!>             @������������������������       �      P�             �?]       `                 �)Ì?���W�=	             "@^       _                 ���?�w���=              @������������������������       �                     �?������������������������       �      �:             �?a       b                 �#�?h�A�R�=             @������������������������       �r��Qjw�=             @������������������������       ��煅���=             @�t�bh�hhK ��h��R�(KKcKK��h �B  '�����>�C���>�Į�N ��.��[~�?� ����>���� ?������?�@���[̿r�� j?����xX忤�`!aW�0UJ�&1? ć`��F?p#E�X�?�����Y�?��;�U$?]}�[X�?Ak�ڽ�?U����龅,�K�.�Z����#�2�Rn����w&.��r�q�[%?�k��Q�?��-!�W��f	�+P�>��VH�.?s���&X�?��k.;W�n,>dG�׾�Z�빿C[�A�?a��k0+?��AՑ�!?Uun�N9?U����cD?+�`\�Y�?��L�HX�? Pæ��#?�qgʺU�?;8�3W�?9s��:��>`���fW���4?B
 �OֿP��@�?����3@?ڵ�Y0x0? ک$QA?wj�uX�?���l�W�?҄�[����V_#YU忌n^=�U忟BT�[]�?D�c�W��'��	�%�
v~��*��e�N�	�0�� �.��P$�U��cW�j����Ǿc�>�U�?����U��W�#��2�h���t8�ϻ��ܿ'���dX��k�*����Z>�er?�d��W�׃�c�*? �ӽ64?�b��UW�?._�լV�?�*&uiU忢�r���>|}����¹�ߛ����rV忈S�]�����z|U�?�Z�2�U�����V忝��Ƈ2?�� ��?��g4?:���J�?��$p�U�x烘Y�?��Ac<�~ц�������ަU�i����U��ˡ�M�㾤�P4\U忦��kpU忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KKh�hhK ��h��R�(KKK��h��Bh                          @@�?V��z�+c>�           �}@                        ��E�?Z�yfH>�            �l@                        ��;�?}����F>�            �l@                        �윳?;�Z�D>�            @l@                        �$I�?@yP��lB>�             l@                        H?�AA�a>             @������������������������       ��ć�zb	>             @������������������������       �                     �?	       
                 ����?Ӱ���@>�            �k@������������������������       ��J�>T)?>�             j@������������������������       ��B�f)P>             (@                           �? �}WƅG>              @������������������������       �                     �?������������������������       �                     �?                       P5y�?@��0��!>              @������������������������       �                     �?������������������������       �                     �?������������������������       �      ��             �?       0                 ��0}?���ABo>�            `n@       !                 ����?ܥ�'Ou>\             W@                         J�N?sB�%�sz>
             $@                         �u��?p2���y>             @������������������������       �                     �?                        �_	�?�X��E*C>             @������������������������       � zka!�>             @������������������������       �      h�             �?                        Pav?�B��fR>             @                        �ߦ�?n���7>              @������������������������       �                     �?������������������������       �      �:             �?                         ��?r?�}�0��'>             @������������������������       �                     �?������������������������       � |�й�=              @"       )                 �*/�?5_X�6r>R            �T@#       &                  漸?�dJ�Fd>             @$       %                    �?��zLo-<>              @������������������������       �                     �?������������������������       �      �             �?'       (                 H��? ���
>              @������������������������       �                     �?������������������������       �      `;             �?*       -                 �v�?z�{
]�p>N            �S@+       ,                  ��?�:��)v>#            �A@������������������������       ���r��Q>             2@������������������������       �u*��>             1@.       /                 x��?^Ʒ�&d>+            �E@������������������������       ��.���g>             @������������������������       ��ʂp�`>'            �C@1       <                 �D�����E1g>�            �b@2       9                  �{��?r�p��K>&             C@3       6                   s��?���oF>$             B@4       5                 P�?�|ڠ��>             (@������������������������       ��
p��l>
             $@������������������������       � �i&8�=              @7       8                 �1��?��l���I>             8@������������������������       �z���=>             0@������������������������       � 7�{>�?>              @:       ;                 ����?��t?<K>              @������������������������       �                     �?������������������������       �      ;             �?=       D                 �0;B?���D�k>q            @\@>       A                 ��ߢ?��뙼�|>	             "@?       @                 �d:�?��z֐1>             @������������������������       �Д�S*�=             @������������������������       �                     �?B       C                  ���?\��Pd�t>             @������������������������       �@����&I>              @������������������������       ��LW��`>             @E       H                 ��C?�i^3p%g>h             Z@F       G                 !C�?  �]�Ղ=              @������������������������       �                     �?������������������������       �      @;             �?I       J                  �߄? �՚je>f            �Y@������������������������       ��x��lu>             @������������������������       �뢼�c>c            �X@�t�bh�hhK ��h��R�(KKKKK��h �BX  �6�e�>�X���g
�y��6OD>�v���g��̥��G �^��4�U��V'?�W�,Z�Yy��W�ݱ¿FC$��  7�
�2?�!<�rW�?���#NV�?P��n:�y���IW�=���W�<�zRW�?_�g&�>d���?:�����5?�wkC��A?�hb�U� �s�`F?9w��[Y�?�͜6X�?�ԓ�"�?�������h1��U��~���U�?�*�n,?8a�V�?惱��V�?���8r?~�F��5�6��?#�q����V��=�j�U�pW�'�@����[X�={��W� ���jT?�z|��� ?���2W�?s�����?'���Bξe���W�?���_$qĿ2C�e�ھ�߱2��\������D��o���:�1�U忘f�U�?�60��&���KV��AjP�V� ���d0#?� .��V�?XU���U�?�[���>��>Ӕs,?T�]=ad�!	�xU��ϡ`CV�fuwܾ<?�=�`Y�?���`W�?��rg�̾���v�=��ݽ
�W忌�I��W志Szy���>>�2'��Cl�M�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KEh�hhK ��h��R�(KKE��h��B                           �`>R?tV�k>�           �}@                        �@�F?v�B3�Xo>             7@                        h�[�>�8���c_>	             "@������������������������       �                     �?                        <�#�?�]� �Q>              @       	                 �I?i~OdH>             @                       @OTZ<?$�֝�'>             @������������������������       �                     �?������������������������       �pi�܍�=             @
                         `���?`����d>             @������������������������       � �Es���=              @������������������������       �                     �?������������������������       �       �             �?                         �3��?�M�Q3Ik>             ,@                         ����?�u��ݜB>             @                         �u��? 
a�r�=             @������������������������       �                     �?                        DWs�? RW"��=              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                        �3M?�9٣f>
             $@                        @�S�? ����N>             @������������������������       �                     �?                        $��?��q�1>              @������������������������       �                     �?������������������������       �                     �?                        �<��>�oh��T>             @������������������������       �                     �?                        N��S?��(>             @������������������������       ��,��b�=             @������������������������       � 9�� �=              @!       4                 �j�a?W+�Rl�k>�           |@"       1                 0��?��Ӧ�v>             3@#       *                  �9��?��[@Ip>             1@$       '                 `ڡ?�<�)�hc>	             "@%       &                 ��^^?e.�V>             @������������������������       �࿛I->             @������������������������       �ƛ�*F>             @(       )                 �l.�?��N���C>              @������������������������       �                     �?������������������������       �       ;             �?+       .                  �~��?�Ϲ��p>              @,       -                  �a�?��oA;V>              @������������������������       �                     �?������������������������       �                     �?/       0                  `���?�7��QAE>             @������������������������       �2����2>             @������������������������       �N�3�#>             @2       3                        YF�-�=              @������������������������       �                     �?������������������������       �                     �?5       6                 ���a?yq �j>�           �z@������������������������       �                     �?7       >                   E(�?~��>�i>�           �z@8       ;                 �R�*?�_�(�f>m            @[@9       :                    �?�<X�dq>6             K@������������������������       �4�<B:h>             :@������������������������       ���l@�s>             <@<       =                 @F�đ�‏J>7            �K@������������������������       ���2�N3J>             :@������������������������       ��U�S��D>             =@?       B                 ��Ԛ?�&����j>@            t@@       A                 �q�?�^ک�s>�            �`@������������������������       ��k�ׂ=p>~            �_@������������������������       ��ɉ����>              @C       D                 `���?��ڙK'a>�            @g@������������������������       ��Kg��q>             :@������������������������       �$u�RY>�             d@�t�bh�hhK ��h��R�(KKEKK��h �B(  ��[w�^׾�'�,�V��8�?�W/�W�? 
@��o�>�h��?|��o�* �!̻��U�?�����U快j���%?s�RV�?7T��V�?ގ`3eV�'F��w)�q,&o��>�w��J�TM�U忁Yd���������U��>�?}U��BQV�?k�^,fT2���@�K��\TW�e{vC�0՚��X��7��9X忲��I'����X�Ei�R �dW?��U�;\J�iV�'����x���
��[L?�V�~'t#?U�)Cq�?������?d�NYV忬��V���?  0{3?
�A�rW�?�eJ^fV�?�3	r�1? �w<�9E?�,X�?xD
�Y�?�G�Ǜ#?-)#`�V�?��X���?X[xNX;�԰U`�W�x"�~�W忰SdCKվ�!�uY志ֵ�˾����3	 ?i�5�?7u�r���?^=���?�}������$�����RB���^�?rY�5��х������￿H�ߕV�߿�Xx��U�>�5j�SM�?�)�� {���t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KEh�hhK ��h��R�(KKE��h��B                           �`>R?m-N�r>�           �}@                        �@�F?���T+%p>             7@                        h�[�>fF��1�b>	             "@������������������������       �                     �?                        <�#�?<o>�4�W>              @       	                 �I?���c�PG>             @                        �~�?�֛J(>             @������������������������       �                     �?������������������������       � K��g��=             @
                        �;�?��?��X>             @������������������������       � ����Q�=              @������������������������       �       �             �?������������������������       �                     �?                         �3��?(��~(k>             ,@                         ����?/1��\@>             @                        �=��? �\G�!�=             @                       `��>�? 
�����=              @������������������������       �                     �?������������������������       �                     �?������������������������       �      к             �?������������������������       �                     �?                        �3M?�v�X��e>
             $@                        Y>t?�Z�h�gP>             @������������������������       �                     �?                        ���J?�bT��2>              @������������������������       �                     �?������������������������       �      P�             �?                        0_Q? @v:	T>             @                         ����?0����R)>             @������������������������       � �����=              @������������������������       �x��\d,>             @������������������������       �                     �?!       4                 �j�a?�O�r>�           |@"       1                 0��?d��F�u>             3@#       *                  �9��?�cyjun>             1@$       '                 ���p?��0�t�a>	             "@%       &                 ��^^?u)v}��T>             @������������������������       ����,>             @������������������������       �jv��̷@>              @(       )                  |�Z?@
����O>             @������������������������       �B�M���7>             @������������������������       �                     �?+       .                  �~��?*��T'n>              @,       -                ��r�?�`��jT>              @������������������������       �                     �?������������������������       �      h;             �?/       0                  `���?�X�a?�A>             @������������������������       ���p�1>             @������������������������       �H�-	/q>             @2       3                 ��[? ��	���=              @������������������������       �                     �?������������������������       �      @�             �?5       6                 ���a?�'}~?�q>�           �z@������������������������       �                     �?7       >                 ���p?V����lq>�           �z@8       ;                 ��"?8YҔ2u>"             A@9       :                  �P��?nn]�%��>	             "@������������������������       �v�@y>             @������������������������       �ԡ���x>             @<       =                 �$?�T(�a>             9@������������������������       �                     �?������������������������       �{{ �*d[>             8@?       B                 ��a,?�˰'�p>�           �x@@       A                 ��j�?_%���Js>�             f@������������������������       ��0FS�fn>7            �K@������������������������       �����Vt>y            @^@C       D                 @��8?~TdD"�m>�            `k@������������������������       �/������>             2@������������������������       �H�&=�h>�             i@�t�bh�hhK ��h��R�(KKEKK��h �B(  !�[L&4�>Ufj��O?��F.���v�m�W��LPS��߾��37.
�5j2��� ?9���U�}���U�?ѹ�B�$���!V�ٴ�\V�zu`�V�?+�k���*?��-��ﾫj�N`q? �rte ?s�ăU�?/�Y~U�?&�n�U�?����=V�f<ct%3? P6�S0A?�]�WW�? ����C?��xDX�?�����X�?n*��<)? `�v�p"?|�6vV�?��+m�U�?����X�?rʗ��ξ8O���W��%#���#���#���}� p�?JQ��ZV�?g�Wim��>/���'�O�v=V�`̧PKW忴�����1��-p�k�D���P	�Y�[60�X�Ag�>�f#�n�o��V���X�U� �_/%�;?�	�h�W�?"7��W�?_\L��ot>g��Y�?ҸƢp����B���?�!��5?�_�qi	ۿ0|^*Y�?mȆ!���X|'��W忑�VY�D�?^3R��ྰy4��S��ֲ���տ�������	��Z�>���W9�? �o�J�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KMh�hhK ��h��R�(KKM��h��B�         "                 �6Sz?w��R>�           �}@                          p��?�gi��R>           �w@                        �lw?G�ZXR>[           �u@                        �ݤv?|�q�Q>V           `u@                        pA7�?��[�l�Q>U           Pu@                        �S'�?�1V��Q>N           �t@������������������������       ��܀���P>=           �s@������������������������       ��aEY>             1@	       
                  ���?{Gr�$@>             @������������������������       �h�z�(>             @������������������������       �      0;             �?������������������������       �     ���             �?                        �q�?�<#�o�V>             @                           �?�?<S�>>             @������������������������       �                     �?                       ����?�s#<��>             @������������������������       ��{S(�	�=              @������������������������       �                     �?������������������������       �                     �?       !                 ���?�C�~XKR>$             B@                        P�bf?����nG>#            �A@                        �r>�?�����.+>             6@                        �t�?-�&>             &@������������������������       �n=��#��=             @������������������������       �x?'i�O>             @                         @�9�?�mx�>             &@������������������������       �H�v��	>             @������������������������       �F<�u��=              @                       �Ck�`?�͡)�FR>             *@������������������������       �                     �?                         �b'�?,R��/8>             (@������������������������       ���U���0>             @������������������������       ��6q/G&>             @������������������������       �      P�             �?#       >                 8�C�?��˨�Q>Y            @V@$       1                 �;�?�.��	�E>9            �L@%       ,                  �Mm�?��U,d|6>             =@&       )                 ����?�Rݺ��6>             7@'       (                  A�?���h�H>             @������������������������       ����A&>             @������������������������       � ��n�l>              @*       +                  �6�?�c�:��$>             2@������������������������       ����A.>              @������������������������       �(o5�5 >             0@-       .                 0��?��ه3;
>             @������������������������       �                     �?/       0                 ����?�LƑ l�=             @������������������������       ��z���=              @������������������������       � ����=             @2       7                 pW��?H�I���K>             <@3       4                  �i�?��/ٞmm>             @������������������������       �                     �?5       6                 P���?`g�ĥ��=             @������������������������       �                     �?������������������������       � ���zZ=              @8       ;                 ���?G�q�*,>             8@9       :                 �O[�?oL|{Ae�=             &@������������������������       ��^�`l�=             @������������������������       ������=             @<       =                 ��^�?ȅepX�5>             *@������������������������       �                     �?������������������������       �YY�^��%>             (@?       @                 ����?�@��ʱZ>              @@������������������������       �                     �?A       F                 �C�? x���.>             ?@B       E                 pl�?D/�m��>             @C       D                   +Y�?���;	�=              @������������������������       �                     �?������������������������       �      �             �?������������������������       �       �             �?G       J                 x�׀?����,>             <@H       I                 <���?��([��@>             @������������������������       �                     �?������������������������       �{N�Uy&�=             @K       L                 x��?o�|�� >             7@������������������������       �ΓM%��=             0@������������������������       �P�9R2>             @�t�bh�hhK ��h��R�(KKMKK��h �Bh  �D���>��w��ƾ�ɷ��0d��پ���7޾�{���U�~�9��G,4p��ݿ�p��?�*mU��?�����V�?B(ư W�?���"�P���u�1F��U�?��u�~� ���8��U�Ko6�>V�Mݲ�xW�]��	?��w��?	�X>4`˾��Ε�����dSlU�y,��U�t��i?��$�U�?H$b�uU�?U�(�?�A�W�?�0i�?5V�?;QF,x�?��2X�?�%�N�R?K�E��?X���G?�i�t�D?3�[d3�%?�TY$�U�?t����V�?����e)?���{DV�?L�L��U�?�j�}��?�cD��U�?�L�h�5�>�=�bU�?�q�ԄU�?�{NM���>���^��a��
X�U�+�u?y�loxU�?�iߢ�U�?U%��s�?F�Er���>_��8jU�?�W���U�?��ֻ>�?���V�?��ֿ�U�?HC�����v����Y�a�E�ƌ�>��>c�? `y�?>\QŪU�?=�JU�?�o7��U�?��	V�s�>��������{V�z���lU�?�o����>D�b��U�?s�>3[JԿ�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kmh�hhK ��h��R�(KKm��h��B�         4                 )DW?�k�!��`>�           �}@                        ���p?�oV��S>b            �X@                        �X�"?��%zO>-            �F@                        �j�a?�
j�P>!            �@@                        �$?Z?�7��#k9>             7@                         �3��?T����r3>             0@������������������������       ��C��C&>              @������������������������       �1@��8/>              @	       
                    �?��$�:>             @������������������������       ���؎�H!>             @������������������������       �      0�             �?                         Ӳ?��6z��X>
             $@                         ����?F/���Y>             @������������������������       �D�F��/E>             @������������������������       �                     �?                         �P�?p~h��L >             @������������������������       �P�K�@>              @������������������������       �   ���<              @                        �$?d� ��j8>             (@                         ���?Q�39P>              @������������������������       �                     �?������������������������       �       �             �?                        0��o??r�(2>
             $@                        pD`n?4���>              @������������������������       �$W�Zu/�=             @������������������������       ���4����=              @                         ��?���	&	>              @������������������������       �                     �?������������������������       �      �             �?       %                 P��{?�vF��T>5            �J@       $                 ��{?A�T�SC>             2@        #                 ���z?�pJ<q;>             1@!       "                 @fQ?�l�qvD7>             0@������������������������       �@$);�3>             &@������������������������       ����p�">             @������������������������       �     �S�             �?������������������������       �      P;             �?&       -                  ���?��KV>#            �A@'       *                 ��<�?����K>             >@(       )                 ��$?�8o9�O>             .@������������������������       �V���ڊ4>             @������������������������       �4����D>              @+       ,                 �-�?4%�d�<6>             .@������������������������       �� l`�I1>             ,@������������������������       �      ;             �?.       1                 x�R?���)`>             @/       0                 ��B4?��(g-4>             @������������������������       �P%�3�=              @������������������������       �       �             �?2       3                 �b'�?���r~0>              @������������������������       �                     �?������������������������       �      @�             �?5       P                 0S�r?���QZ~b>v           `w@6       C                 0���?��f�c>�             d@7       >                 P��?�[�ȭ�h>Q            @T@8       ;                  �G?�?���ݗBg>L             S@9       :                 ����?J����/e>B            �P@������������������������       �<�p�ib>>             O@������������������������       ��Q��m>             @<       =                 ؿk?O���bi>
             $@������������������������       �                     �?������������������������       �$�R�e>	             "@?       @                 ��7�?�'��w`>             @������������������������       �                     �?A       B                 �m��?0r(!�EE>             @������������������������       �                     �?������������������������       ��� M�$>             @D       K                 PĚ?'�/^V>P             T@E       H                 �5�?C{$*3d>             *@F       G                 p�3G?�N8��+c>             @������������������������       �x����)_>             @������������������������       �`v_bZ�=>              @I       J                 �؉�?�59���'>             @������������������������       �.t���>             @������������������������       �       �             �?L       M                 0N��?��_�L>C            �P@������������������������       �                     �?N       O                  0C�?bN&��<F>B            �P@������������������������       �                     �?������������������������       �v+@�?�C>A            @P@Q       ^                 �&�?��3��a>�            �j@R       Y                 ���6?�qg6i�c>g            �Y@S       V                     �?�E]n�.d>-            �F@T       U                 ���?���A	zU>              @������������������������       �                     �?������������������������       �      1;             �?W       X                 @ܒz?4.J�a>+            �E@������������������������       �3E�-�tC>
             $@������������������������       �4KL�a>!            �@@Z       [                 j:?�\�c�`>:             M@������������������������       �                     �?\       ]                  �_�?�΍�>cZ>9            �L@������������������������       �,���o9>'            �C@������������������������       ��x�'�n>             2@_       f                 �c��?�ɣLg�\>n            �[@`       c                 ����?���ʏR>             @a       b                 ��-�? `�>��>              @������������������������       �                     �?������������������������       �      0;             �?d       e                 P��?���E;>              @������������������������       �                     �?������������������������       �      �:             �?g       j                 �Y8�?%�F��[>j            �Z@h       i                 0?�����v>             @������������������������       ��A��ea>              @������������������������       ���&�[+>             @k       l                 �H�9?�>
�.�V>e            @Y@������������������������       ��w���q>             9@������������������������       �؏�W��2>L             S@�t�bh�hhK ��h��R�(KKmKK��h �Bh  ��N?��¾��m�:�>��MaXFﾜ�U�t��=����>�W�L���Q�Ͷ��?�����{����$
?m�����?4��#}V�?9ϯgt�"�o/�ig�+���0]��w� JX忢�"����<�c�?����U�'6�@N�? 
Z��#?J�q@�V�?�봮zU�?��h�d�?rB�^C�>�G?�U�?�D��oU� @��H?�A\V�?W�&��U�?�{@b�?��ґ� ?�igH��? ! ?��V�?`]�NdV�?�b�wU�4�EW�?�.7N ?��৾$�>�jP�xW�G�\#o�?��G0�\sΘ��?��ۻ���?�껒�U�3�0�f+?UIz�u?1���U�?T��HV�? \�g�:?�WL�5W�?��<P�W�?�*��%#�O@����4_VR�������?̢%���s̰ѿK@��3��?"����i*���x�8X��kY�+W俾� �JC4�C��_U�ڱp��49��D�RIX忷�Y�0W�E
Y���>nv�;��"?%9�D�O1?��7K5W�?�����W�?]����>�1��U�|"��U�?N$oT��2g��W忮F�$��Hy��V�?���&�ǿLu08�M�>ұQ�O�?�Ts`�? }�S;�,�F��`LW���
��U��R>.;O ?;����+�q�n�?8�O������G�X��������>�Up�ۿݜ�r�?�?߬ڥ������*�1M�q�$5���AW�zu$S�V忘E��
4����@V忨�UbU�|�_����C��&?�M�iX�?���O�U���`Y(������tտ��:z�y���t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K]h�hhK ��h��R�(KK]��h��BX         4                 �SpR?�v�g�f>�           �}@                        �U����$���[>S            �T@                         W��?�K�EA�c>"             A@                        ��??y\j闋Y>             9@                         .:q?���mL�L>             6@                         e	a?r)�zB�M>             0@������������������������       ��j��n@>             (@������������������������       ��aE�`&>             @	       
                 �Q�?���n*">             @������������������������       �`�r	�
>             @������������������������       �       �             �?                        艝�?�X���e>             @������������������������       �                     �?                        HeT�? ��Xv�@>              @������������������������       �                     �?������������������������       �      0�             �?                        ��ߗ?~G)/�Zd>	             "@                         `���?�@!�(yN>             @������������������������       �                     �?                        k�_M? �Y*)�B>             @������������������������       �                     �?������������������������       � bݣ?� >             @                           �?����L>             @                         p�{�?�7K�ĝ >              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �             �?       +                 ����?�q"�[�F>1            �H@       $                 ��=�?]nf���@>,             F@       !                 ��B?~�4>             0@                         `�լ?Fp[ֲ,>             (@������������������������       ��lY���=             &@������������������������       �                     �?"       #                 ��L�>�}��N>             @������������������������       �                     �?������������������������       ��TOc��=             @%       (                  �"�?��n�gm<>             <@&       '                 ��37?���U�\0>              @������������������������       �l���>             @������������������������       ���x2��>             @)       *                 ��2?T��S8>             4@������������������������       �G\�6_:>             (@������������������������       ��<2:*C>              @,       /                 ��j�?����P�M>             @-       .                 Ћ��?��G$&��=              @������������������������       �                     �?������������������������       �       ;             �?0       3                 @iD?V�a�֐D>             @1       2                ��T�? �,Km��=              @������������������������       �                     �?������������������������       �      �             �?������������������������       �                     �?5       N                 ��_i?R6wxp�h>�           Px@6       ?                  �~��?��_h�[P>&             C@7       >                 P��?��N�@�E>             4@8       ;                 ��V?�t��FvB>             3@9       :                 �9>?G}��~J>              @������������������������       ��{��F$D>             @������������������������       �       ;             �?<       =                 b©�?��:,dT>             &@������������������������       �pxh@�>             @������������������������       ���| >             @������������������������       �      0;             �?@       G                 0j:�?���4�P>             2@A       D                 P�a?Jl\�<R>
             $@B       C                 �w�_?�9�B�PN>             @������������������������       �`k��e�:>             @������������������������       ��������=             @E       F                  `��?@E�R�>             @������������������������       � @����=              @������������������������       � ��7���=              @H       K                  `��?��]��>              @I       J                 ��ǻ?��3S>             @������������������������       ��(聕�=              @������������������������       �@�Ӄ�H�=              @L       M                  ��?��V��=             @������������������������       �                     �?������������������������       �T�!�î=             @O       P                  ��i?d��IKIj>_           �u@������������������������       �                     �?Q       X                 �-�~?p�<�&j>^           �u@R       U                 ���{?-|�Õ^>2             I@S       T                  ���?
C�z�T>0             H@������������������������       ��C�(��N>&             C@������������������������       �Ȁ�~�[>
             $@V       W                 ��?��l�	d>              @������������������������       �                     �?������������������������       �      P�             �?Y       Z                 pk?k?ɪ�&�k>,           �r@������������������������       �                     �?[       \                 �;�?�R��Kbk>+           �r@������������������������       ��[�GPq>             7@������������������������       ��w���^j>           @q@�t�bh�hhK ��h��R�(KK]KK��h �B�  p�W�N���>�$��>�F忤�?v|��?�����>���@F	?��
�ΐ�7��n|V�?'�X��?��U�	��.V� p�Z�#2?�2��dU�? ܩ��:?_�$0X�?��W�?�ٹm.�1? ��@�8?��0dV�?�ў��<;?���l�V�?7~5�W�?��{�L0
? 8c$G� ?�ow2�U�?�}�5EV�?�À��U�
�x���ќ��@���H���>ޢ}������t�U��4HNOV�? �7�s3?]}�+V�?����U�?����kf�S��;�l��j���U忔=ܶU�?�lv����P�sh��R���+V�8I�L�? �d��?-?آ��V�?fx+�uV�?4��aF?ңQ����FRtzU�HG6�U����OV�?���9��ھ|T�+}e�����r ��&p�䙽�� ��-�>���b$��C:NacV�?�M@�����Ɂ�U忩�ҮU��~�:V�?�ˮ�I� ���;�Z)�XuM=j��A�b��V忈�q{U忇��3&�3�Q x��V��h�/W��F�ݾ�B_P�`��)�If�U���x��U�c�أ�1�Կ
�U�2u*;bU���閮>1O�WZW�?v�.�g�������	?�p&G���>5H3��?/(t;�? ����5@?C1��V�?�o̯Y�?�N�\�l���9�X����Iܾ������?ꚲ�簿�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K[h�hhK ��h��R�(KK[��h��B�         6                 pY7e?�5T5>5K>�           �}@                        @E��?�]��@�L>h           �v@                        `ӣ�?�0��[�J>(           �r@                        �!�?�;�L��F>�            �o@                        ���?IMr�ȠB>�            �n@                        ��?�bߍA>�            �l@������������������������       �N8��h6>�            `j@������������������������       �MA�{oc>             2@	       
                 �7?���'~N>             1@������������������������       ��UF�ca>              @������������������������       �����@>             .@                        h��1?{0��]�o>             @                        8�2�?��Gx�^L>             @������������������������       � T����>              @������������������������       ���/��=             @������������������������       �                     �?                        �!�?��H_HV>,             F@                        ��h�?�$�]P>#            �A@                         �E�?�qG>"             A@������������������������       �o��(��7>             ;@������������������������       �/��GY>             @������������������������       �      l;             �?                        �\��?�1���[>	             "@                           �?P�۝RB>              @������������������������       �                     �?������������������������       �                     �?                        p5W�?��ܭ�&>             @������������������������       ��wFx�t>             @������������������������       ��1�w�+>              @       -                 |�L?��F}w'S>@             P@       &                 �v�?Oe�V>!            �@@        #                   +Y�?�
: ߘ`>              @!       "                  y��?4���ĽV>             @������������������������       �@�5��>             @������������������������       ����/�0>              @$       %                 `���?8�����=             @������������������������       ����"~��=              @������������������������       �      к             �?'       *                 P�8�?���xA>             9@(       )                  P�J�?��tk!8>             @������������������������       �F�V�LZ>             @������������������������       �                     �?+       ,                  ���?�j-�;>             5@������������������������       �                     �?������������������������       �&q�g+>             4@.       /                  e0�?��*�F>             ?@������������������������       �                     �?0       3                   +Y�?P����@>             >@1       2                 ��ލ?	/��&2>             5@������������������������       �8�H �0/>             @������������������������       �Rx�}p�#>             0@4       5                   B�?�B��BC>	             "@������������������������       �                     �?������������������������       �� t��N2>              @7       D                 p�m?���'�D>p             \@8       C                 ����?��K��i>              @9       >                 X�E�?�4���[>             @:       =                  pS�?���p��>             @;       <                 �.�?Ht�!m�=              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �             �??       B                 pU�l? ��4|�H>             @@       A                 �m�? \$�s�>             @������������������������       �                     �?������������������������       � ��b��=              @������������������������       �                     �?������������������������       �      X�             �?E       L                 p�,p?N�ݞ�v9>h             Z@F       I                 ����?h�fzU>             @G       H                 `���?�P J\@>              @������������������������       �                     �?������������������������       �                     �?J       K                 p~�?��r ��=              @������������������������       �                     �?������������������������       �                     �?M       T                   �?Tz��85>d             Y@N       Q                 �Ys�?�e�ەB/>@             P@O       P                  ���?2�H��  >/            �G@������������������������       �dI��_>.             G@������������������������       �      0;             �?R       S                 @�	�?o��&N�?>             1@������������������������       �N�]lO�T>             @������������������������       ��Y�O�a>             *@U       X                 ����?�)�J��;>$             B@V       W                 h�؝?7�-���`>              @������������������������       �                     �?������������������������       �                     �?Y       Z                 �ܳ?4�"Aw>"             A@������������������������       ����,>             @������������������������       �C���*�>             =@�t�bh�hhK ��h��R�(KK[KK��h �B�  OG2J[�>��nmƾ_N�K���+��«��Q�|O?پcuYI����T�'TĿ�j���z�?�;c��Q�Q_W�d�;��ۿ�*>H��&?����E�?��ބV�?�5��yU�QX���X�?q�\�\���:ߎ���������L|(� ۚ�
�ῲ6���W�'z���? (Ku��6?���V�?�Kc{�W�?�S[��ݾq�`*�U� 0��q�?th"�>Em0׵�? �B��,? ��*d5?I?<V�?o)�X�?Uk]T�?-ʗu�U�?w>�|qU�?��f��>e�1�<�����S�U����sV忄첑�?T*���V�?��5�2Q�?qT,�o��Cs�U�V�?�M3�& �ց(Sd7��et�5V� �"���{��R�?���V�?UY���@�?p1� ��>�+�N ?�����'?�-ݎ�;�> �"�`?N�B�U�?C6��U�??x�U� V���3? P.Z��/?���UV�?r����V�?݊*�W�?�m���V�ĪZ\h2�>�������U�Vs,�Ÿ���V忍I>�
V� @Gy�e?���U�?0�UzU�?���[��>*$�
��>��0*2C?�E�Cu��?�sDV�?�w5�n0�� $�5�ܿl����U�?Na���A=�/�'8ۃ�U�k�Bl�W�a��>��4�ֿ�b���?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KAh�hhK ��h��R�(KKA��h��B8         @                  @���?,Y�ڐP>�           �}@       !                  ����?�S��zP>�           p}@                        ����?n��3�JU>           �q@                        ����?��و�d;>g            �Y@                        @F�O7}2->9            �L@                        ���L?	�����%>$             B@������������������������       ��=�6��%>             6@������������������������       ����ԙ�>             ,@	       
                 P�r?�p,+�0>             5@������������������������       ��f)�9>             *@������������������������       �6>��I7>              @                        `��?���#�B>.             G@                        �-�?�E~�J@>             @������������������������       �8<Ĩ��>              @������������������������       �                     �?                        p#��?PVb�ӥ?>+            �E@������������������������       �������E>             *@������������������������       ��@F �23>             >@                         �~��?�z^��\>�             g@                         (V�?�Fn�bP>v            �]@                         ��~�?*.t+�#P>r            �\@������������������������       �                     �?������������������������       �փ�$w�O>q            @\@                        �h��?��ވJ|3>             @������������������������       �����=              @������������������������       �Lo7U�>              @                          �P�?ᥪ�h>B            �P@                           �?�P�f�>             &@������������������������       �� {�%�>             @������������������������       �O��g�=>             @                         p���?��5�*�V>7            �K@������������������������       �����#�Z>             8@������������������������       ��(��dP>             ?@"       1                 �y����'�-�yA>�             g@#       *                 ���y?<�-��M>C            �P@$       '                 ����?�b�+BG>/            �G@%       &                   +Y�?��!�x�G>             <@������������������������       ���M��Z.>             0@������������������������       ����f�Q>             (@(       )                 ���?�z8�:>             3@������������������������       ��M�N�>>              @������������������������       �ܻ��>             1@+       .                  Ff�?z��CR>             4@,       -                 (��?.�݂�H>             ,@������������������������       �zB��~�>>             &@������������������������       �q`s�}�0>             @/       0                 ��}�?�&k�9-;>             @������������������������       �                     �?������������������������       �\���gN>             @2       9                 �f1�?�ԑl��4>u            @]@3       6                 `�w?D|�E�->             5@4       5                 `@�_?��]>Q�=
             $@������������������������       �8�L���=              @������������������������       ���
o!P�=              @7       8                 �|c?���U�s3>             &@������������������������       ��%mF�T>             @������������������������       �`i=iW84>             @:       =                  p�:?/��/�3>`             X@;       <                 P�$�?�#Fh��S>             @������������������������       �t��I�J>              @������������������������       �                     �?>       ?                 ����?K =�р->]            @W@������������������������       �$+��>/            �G@������������������������       �z7y1j�5>.             G@������������������������       �     �û             �?�t�bh�hhK ��h��R�(KKAKK��h �B  �t��]>�%]�����
�H,�>�]X�����v,`�>�t8�[ݾ%�����?���~�U�4o��Y?]�?m�#�?�$\��?n���a�U���lA?6ӶL�U�?���~V�?̴��S�׋������I��%�߿[Hy���>	A��7�>0p��!�>T�穛V�?	�Z��f�?o��`� �����aV�ϼ@��U忁��ԑ>?�q�J�%?�
S���?)��I���y��X�>N\�� ��?*/H���z��d:�m�$�0�������y	��E
ب��UG���W�cj���g��>�S-֖V�?��֑�U�Љ���T�>�#��?�1gg",�?�pG��ῌ� q���[m�V�����U���.HGž'�$��?!�5��>1�sU�?�ׁ�oU忺( �M�?�ڰ�U�?�ʣ�BV�?9�;~�龻ք7�d$�X<��U�Rg��1W���mO��߾y����U�Y�u�?�#��V�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KUh�hhK ��h��R�(KKU��h��B�         &                 �C�?O	��U>�           �}@                        P˦�?���{��W>x           �w@                        0�P�? ���W>V           `u@                        ��ذ?�%&�)W>S           0u@                        ��n�?4��\(R>=           �s@                        ��{�?��:�Q>           �p@������������������������       �Cs}DQ>�            `k@������������������������       ����eu�M>3            �I@	       
                 Z��?NM��V>/            �G@������������������������       �                     �?������������������������       � 2���R>.             G@                        ���?��|B��v>             6@������������������������       �                     �?                        ��^o?�V�p�K>             5@������������������������       � ��6�Ԕ=             @������������������������       �v4��vA>             2@                       ��ח?`a�ҳM>             @                        �/�? J��<a�=              @������������������������       �                     �?������������������������       �                     �?������������������������       �      P�             �?                        ȬH�?��BJ>�T>"             A@                         ����?��0Ct�O>             =@������������������������       �                     �?                        PL�? �[?p@F>             <@                        �xȯ?@�Br=I>             0@������������������������       �+����B>             .@������������������������       �      b�             �?                        �ٰ?�!��&�1>             (@������������������������       �                     �?������������������������       ���-��>             &@        %                 '�g�?�Iv�G>             @!       $                 `TF�?�Ee\:A>             @"       #                 ��J�? �Qp�=             @������������������������       �                     �?������������������������       � �18��=              @������������������������       �     `;             �?������������������������       �     �#�             �?'       :                 ���?��ŴGDJ>`             X@(       7                 �и?�O'�bV>             9@)       0                 0��?�3��u3S>             7@*       -                  e�?�Z�e�^2>	             "@+       ,                 `h"�?���m�0>             @������������������������       ��v�T)��=              @������������������������       �0�����>              @.       /                  �g<�?"�dbC�>             @������������������������       � h���,p=              @������������������������       �P���x��=             @1       4                 ��;�?����$�W>             ,@2       3                 lH�?��4�o�>              @������������������������       �                     �?������������������������       �      0�             �?5       6                 `s5�?�M���J>             (@������������������������       �����[0>             @������������������������       ����O>             @8       9                 g<�? h(b��=              @������������������������       �                     �?������������������������       �      0;             �?;       F                 ��? �ÂB>G            �Q@<       A                 @}wL?�o{��`>
             $@=       >                 ���?n���f@Y>             @������������������������       �                     �??       @                 �#e�?� �V�0@>             @������������������������       � :���>              @������������������������       � �����=              @B       E                  ���?(57U�D>             @C       D                 A�Ӛ?�P�8�>             @������������������������       �                     �?������������������������       �@�W*���=             @������������������������       �                     �?G       N                 `L?���<�!0>=            �N@H       K                 Pg�?��	��)>             8@I       J                  �@�?�xe�$�>             5@������������������������       ��Y9�eg>             4@������������������������       �      $;             �?L       M                 ��R=? :�/�>>             @������������������������       ��bd���=              @������������������������       �                     �?O       R                 p��z?D�����0>%            �B@P       Q                 �1Nu?�=ܪ�D>             &@������������������������       ���1��/>
             $@������������������������       �                     �?S       T                  ��?�GQ7�>             :@������������������������       �                     �?������������������������       �k���[�=             9@�t�bh�hhK ��h��R�(KKUKK��h �B�  $_��벾�Ɂ*ڃ׾RMt��B���w3c��ʾ��z��>��uGy߾2T��L>�?ӎ^�ؿL(fRj?�w{�W�?L�;��5�?M�	�~�����eX\��tA����>
�x�SV�pR�'���?����M�1? �||%�(?�~�AV�?K(6�wV�?��>�W�?���׾8���38��=s�W�mG�l8����/��1�1v[V忸9�A,W�,���ĥ��c$��1V�?IU�U忣�H��?%�y�J#?U5�*?YF�RV�?��wV�?���^U�?��sU忳0sl�5�>��<c�
?���-� ?�����h�h����v�c����U�:?^$V��K.��>����U�?J��xU�.7>? ���B�5?���!WW�?͏���V�?+6Obn��>N;��U忥�b�A$�? �f}�2?$1_2�V�?.�uq�V�?�X1�=k�>�p��?�y��*?,V"-�U� �q6�1?{Љ,FW�?�8��UV�?���}c$��K|c��>-�2E�U�?�g��hU�f} J�V���j�0c����r_���:ˊ�쾫������C?Q��U�?�AvĆ �*��U�0YCWV��m���>�1��*c?z��Hb��?Z��V�?ֈ�!�r���U� zgsU忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KSh�hhK ��h��R�(KKS��h��B(         &                 ��K�?ڭ�T6>�           �}@                        ��?��V�?>�             e@                        �\�?����<�>k            �Z@                         �.�?�z�,/�=Y            @V@                         �F�?jFi��=X             V@                        ���@?���"��=S            �T@������������������������       �Z�9)�j�=@             P@������������������������       �fO���1�=             3@	       
                 �Og�?�dOP~�=             @������������������������       �                     �?������������������������       �@4g+��=             @������������������������       �      (�             �?                        `e�?���p�@>             2@                        &yP?�*���K>             @                        ����?�N�)�L>             @������������������������       � ����>             @������������������������       �      -;             �?                        ���{?( �[�>             @������������������������       ���\�o�=              @������������������������       �                     �?                        ��h�>|�:ӥ>             &@                        P\�>�:�(S#>              @������������������������       �                     �?������������������������       �      �             �?                        ��Z?�,�[�=	             "@������������������������       �Jn1%:��=             @������������������������       ������=             @                        ݔ?}!^v��Q>>             O@������������������������       �                     �?                        �$I�?YdU��J>=            �N@������������������������       �                     �?        #                 �3,�?m���DJ><             N@!       "                 �@�?�D�s4T>             <@������������������������       ��"k�d8>             .@������������������������       ������]>             *@$       %                 �mf�?$�]A8>              @@������������������������       ���%b�QU>             @������������������������       ���	g�">             <@'       8                 �7��?C'&��0>/           �r@(       7                 P��?8���"1>�            @o@)       0                 P�$�?DWVg�0>�             o@*       -                 �O�?���M��->�            �i@+       ,                 ��c�?���t'>�            �c@������������������������       �w/�G��#>�            @c@������������������������       ��>�
�Q>              @.       /                 ��E�?����r5>3            �I@������������������������       ���@���5>%            �B@������������������������       ��%�}l4>             ,@1       4                 P^��?j�f�/6>*             E@2       3                   E(�?�. M�4>(             D@������������������������       �K]Lļ>             1@������������������������       ��?yq<>             7@5       6                p�~�?� ��w>              @������������������������       �                     �?������������������������       �      �:             �?������������������������       �      �             �?9       F                 �\��?���Z7�)>5            �J@:       ?                  �˛?{'1�w�'>#            �A@;       <                    �?��n�d�6>             @������������������������       �                     �?=       >                 
�jU?`�C:W�>              @������������������������       �                     �?������������������������       �       �             �?@       C                 �u��?l���y>              @@A       B                 ����?N]�*�?>             0@������������������������       ���! ��>             .@������������������������       �      0;             �?D       E                 ����?���M�>             0@������������������������       �                     �?������������������������       �4(�N�~�=             .@G       L                 �s�?����Z�$>             2@H       K                 �ڡ�?��.4+2>             @I       J                 ���R?Ms�� >             @������������������������       �8�����=             @������������������������       ���*X}�=              @������������������������       �                     �?M       P                 tU�L?g�.��.�=             (@N       O                 ����?�8�7�=              @������������������������       �                     �?������������������������       �                     �?Q       R                 �#�?�,Z:��=
             $@������������������������       ����wb�=             @������������������������       �Ht#u��=             @�t�b��     h�hhK ��h��R�(KKSKK��h �B�  چ&tw�>@�[Tn��> �z����t�G�۾ڊ���׾$���CѾ�B��\U��7��
��΢��� �!X�Y�U����zU忌�/�U������>.wi;�?��̵�n"?��>|V�?���U�5t����>{�# ���n�}�U�?��X}	��LCL���:�iU忬���U�B�S�Bᾍ`��qU�Yh��ڭ�?&\���?6m&:X�?������>�I��V�{������>���?,ܛL=O�?�=��ل�?c�H=��>�Ũؿ���6-��?UR8dE~Ծ����g�㾧����%�D��j��dڏ_��־wX�Rɿ= ���V�?�����O�$��,��-��?�P����>5Ҙ@��>'5��������Cxy�?nP-R���L.�V忮�,��U�̓��aV���u.#�>�3zH-g�> ���b ?���{U�? x�; E&?��-6rV�?ˬS�V�?��RO8�>�P���?��7��q�?C�=9�U�?(���{�>Q��V忎HK��U�?�Ț+IPᾱ��<N�
�=7��$���p��׿�䫞�U��?b]V� �ѷ.&�> `�R�?��s8�U�?Q'U�U�?  9���>�ܼ�\U�?f�jU�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kmh�hhK ��h��R�(KKm��h��B�         8                 0���?�V#��8>�           �}@                        �2*�?�j�8>O           �t@                        p'v�?ʳu��C->�             j@                        й��?����'>�            �h@                        �C
T? �|�i#>d             Y@                        �U�����9�W�>:             M@������������������������       ��H�>             6@������������������������       �})>o>$             B@	       
                 ��??�9'\S%>*             E@������������������������       �(��$>             ;@������������������������       �����N�=             .@                        ��b?��[��"*>c            �X@                         h2a?!����J>             @������������������������       ��	��,X*>             @������������������������       �                     �?                        ��/�?�i�">]            @W@������������������������       ��'�(�B>             @������������������������       ��NL��>V            �U@                        ��*�?"��bKLO>	             "@                        ���N?�]��{�X>             @������������������������       �                     �?                        �*�m?Y3@T��8>              @������������������������       �                     �?������������������������       �                     �?                        �[�?bT�M�>             @                         �a�?����r\�=              @������������������������       �                     �?������������������������       �                     �?                        �Q�?P.B��=             @������������������������       �@��$W��=             @������������������������       �     �к             �?        -                 @C��?�����C>            �_@!       (                 ���u?-��x�G>?            �O@"       %                 pyӂ?�p��/>             1@#       $                 ��ѡ?_�d:��>             .@������������������������       ��8uu�.>             ,@������������������������       �      .�             �?&       '                 �@	�?)�N��RA>              @������������������������       �                     �?������������������������       �     ��             �?)       *                 �m�w?���x�J>.             G@������������������������       �                     �?+       ,                 ֢�?�� ��A>-            �F@������������������������       �)�u�&�=>             8@������������������������       �	}��KXA>             5@.       3                 `�l�?��8�&<>@             P@/       2                 �ڡ�?4AQ8�T>             1@0       1                 �(�?�G"�4?N>             0@������������������������       ���Q:B�N>             @������������������������       ���z$Ћ4>	             "@������������������������       �      d�             �?4       5                 �u�?۷���K>/            �G@������������������������       �                     �?6       7                  ����?v9��i�>.             G@������������������������       ��V!xG�>-            �F@������������������������       �      $�             �?9       T                 ����?��Hˡ�8>�             a@:       G                 �7��?���-��I>             7@;       @                   �G�?}�+n��>             (@<       =                 �vQ?來��+$>             @������������������������       �                     �?>       ?                 �Bk�? ���X|�=              @������������������������       �                     �?������������������������       �      �:             �?A       D                 @2ΐ?����9��=	             "@B       C                    �?Ho��>             @������������������������       ��(�ŋ�=              @������������������������       �                     �?E       F                 ><(�?l�D���=             @������������������������       � �Ǎ�=             @������������������������       � ��/�=             @H       O                 ���?,�Ob%}P>             &@I       L                  �נ?���H)�9>             @J       K                  �x��? ���x�>              @������������������������       �                     �?������������������������       �                     �?M       N                  �9��?`Xq��>              @������������������������       �                     �?������������������������       �      �             �?P       Q                 ���?�S�1>             @������������������������       �                     �?R       S                  (��?ٍ�Z�>             @������������������������       ��ael(��=             @������������������������       �       ;             �?U       ^                 PX�?Auѿ��1>r            �\@V       W                 ����?@E31@�>+            �E@������������������������       �                     �?X       [                 �H9�?P�4�>*             E@Y       Z                 pTF�?ɻC��y>             ,@������������������������       ����֒��=	             "@������������������������       ���E�>             @\       ]                 �:WN?�3�e>             <@������������������������       �oa���>             *@������������������������       ���e���=             .@_       f                 P�o�?@����6>G            �Q@`       c                 `WJ�?D�MF��;>
             $@a       b                 �P�?H��x1>             @������������������������       ��8�4�>             @������������������������       �      ;             �?d       e                 0JW�?�o��J>             @������������������������       �                     �?������������������������       � �"���=              @g       j                 �3e�?�{Z�lJ3>=            �N@h       i                    �?��QF>	             "@������������������������       ����f�>             @������������������������       ��+KZ�B>             @k       l                 �x�?W�j��2(>4             J@������������������������       �: �<�2>             @������������������������       ���CxC">1            �H@�t�bh�hhK ��h��R�(KKmKK��h �Bh  ��1��g��!�jm�վ��Մζ�>`D7�1p�m����>�/�:<�ܾ���	 ڿ�����?3Lk+�j?T&l�l5�?Mz�9���䙲e��Ո�2�?tL [��?�A+}�V�?]�2��B��0NP�r�G���طڿ"i�
�,?3s��>&?XX$TW�?��x�c�?FD�ZU�;C��#V�?}V�7H��  ��a� ?C�BqU�?$h<��U�?X�('��橰AuU�݀�$[U�__&����|<���#����>��h����>��8)���?I����U�x����38PB^V���cU�R+O���I�B�X����Ӵu	�3���b���hH��ſeTg6p�>�q��g�
?�,	Zt ?Ji'<�|�? �Qrֿ"g	IW�?C�{pd� ��tV��[��Qྍ6�&�U忐����U�?�oi���> �W���?O��T$�Ԑ��d���斨V忘A������gxU�0)�qU�d��?-��>J��}����O~k���J��U�UU�m�O�>�v��aU�?:AQ�sU�?DRلe.? \��30? h�d��4?Cv��V�?v��>W�? ��`F*'?�ȁzV�?7��pV�?��'��?����5V�??a�H�>����U�?�����U��ӽ-��>-��\~��i�fV����8=U��mr�u�>\�=��^�?�ru��ٿ��@�5���m!���-�'k�U���䘈�>�ŠV�?]����K ?���
s*�?y7ۙ5V�? �N)Û$?w�S@mV�?�BǑV�?���Js��>��6�b ?�^'�!��%�qZ\��?�v��پo٭� V�R�a"c5E?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kch�hhK ��h��R�(KKc��h��B�         $                   �G�?��k�a?>�           �}@                        @j��?iE�gO3>@             P@                        Pz�?�e�Н,>=            �N@                        0B��?�<N�*>(             D@                        PeT�?����!>             <@                        ��ם?�4*��g>             5@������������������������       �����C�>             3@������������������������       �\�A/�>              @	       
                 @8��?4G����&>             @������������������������       �`��-�>             @������������������������       ��*��>             @                        ����?_�w�/>             (@                        �@�A?1�h|�J>              @������������������������       �9Lח!f>             @������������������������       ���4�zE�=             @                         �G?�?���.5
>             @������������������������       � _7}�=              @������������������������       � �ӑ���=              @                        ����?�b��R�%>             5@                        @�C�?z�F 4
 >             (@                       ��Xv?Lb{(�>              @������������������������       �
�A���=             @������������������������       � �0\��=             @                       �+q%�?@�k��>             @������������������������       ��a��o�=             @������������������������       �      ;             �?                          ��?���v[�>	             "@                        8<o�?�ߙ*>              @������������������������       ��x�9A��=             @������������������������       �      �             �?������������������������       �      �:             �?        #                  p��?*��ޱ�O>             @!       "                 �f�?Ž(X#>              @������������������������       �                     �?������������������������       �     ~�:             �?������������������������       �      0�             �?%       D                  �P��?=/��Q�@>�           �y@&       5                 �U����1��<<>L             S@'       .                 ��Z�?+Ճ�/A>!            �@@(       +                 0��\?���y�">	             "@)       *                 *x?����0��=             @������������������������       � B��lD=              @������������������������       �      �:             �?,       -                   E(�?���п�!>             @������������������������       ��h���>             @������������������������       �      �             �?/       2                 PkԐ?l��CB>             8@0       1                 ��ߓ?�:l��%D>             &@������������������������       �p̒����=             @������������������������       �s
��B>              @3       4                  n��?�mz�,>             *@������������������������       �                     �?������������������������       �Ά�`
M#>             (@6       =                 p'v�?xiE+�/>+            �E@7       :                 (߁C?��05s�#>             6@8       9                 H�x?R�E�@C">             *@������������������������       ����
d�>             (@������������������������       �       �             �?;       <                 �q��?�Ż��O>	             "@������������������������       �=�	���=              @������������������������       �                     �?>       A                 `s5�?��R�1>             5@?       @                 �?�?����֋">             @������������������������       ��a���>             @������������������������       ��6���>              @B       C                 �VS,? �p!'>             0@������������������������       �                     �?������������������������       ����>             .@E       T                  �~��?�W1)�@>L           �t@F       M                 �-�?�1H�ʮM>0             H@G       J                 0I��?<�UE�Q>             ?@H       I                 P���?}%SNM\6>             5@������������������������       ������3>             2@������������������������       ��0�o5�#>             @K       L                 pTF�?X]m�@_>
             $@������������������������       �                     �?������������������������       �H0�z��P>	             "@N       Q                   \��?�p�a8>             1@O       P                 ��j�?0�+u��#>             @������������������������       �`���[>              @������������������������       �      ;             �?R       S                   s��?W%�)�^2>             ,@������������������������       �Z���V&>             (@������������������������       ���jV�8>              @U       \                   �P�?�Z!Q��<>           �q@V       Y                 �D��C�\F�G>             ,@W       X                  �ȗ?o�z��N>             @������������������������       �ې'�ӂ#>             @������������������������       �                     �?Z       [                 @��I?��各�6>              @������������������������       ��/�Im�">             @������������������������       �<�5SS#>             @]       `                  FS?�?>��;>           �p@^       _                 ���?B��G؃3>-            �F@������������������������       ��ӎ�/>,             F@������������������������       �      D�             �?a       b                 ���?��(��<>�             l@������������������������       ���b���B>)            �D@������������������������       ���א�9>�             g@�t�bh�hhK ��h��R�(KKcKK��h �B  �����q>�KEȩ�>��4���>��/�%wҾ1��p:��>=��m�ƾ����D��?)��@�U�8�O�?�̥S�U�?��~��?�>���R[pRB׾�����/߿�5h��U�?�s�Z�[�g��U��"�V�5��ɭ#?��F�7? �T�i?;�ˊU�?_��Z�U�? ��b=?�[�V�?̖ ��U�?/X�C�>�0qQ�ܾL�==*����K�U�_����U�?�q�E�� ?bIG/�?��1��U�?��T�UU忰�6|�V�?��9�Bľ���HE 󾦗��X�M�9a�>��,�S;���P�zU�z�JQ�U������>^�dVTx�?h�7�U�!��QB���R� �h�N��U�Rl�V�I#6@n� �3'L��U�?�|xND��X6E���>O}����꾱)�����kQ���޿IG�a&V忽��H��>�9v=��?� 0W�U�?��	4?  ��q?�S��V�?a��U�?W�&P��>�X�;V�?'ASSR?p�J��˳>�V-8���>n5��|0?��#*��>W\��#��4��+�U�?3���"?i�DY#X�?9`�,�?�_���i뾫�(�*�$�y V�D�+�U快��Y�>�����X�?F6*V��`���Ͼ�bp���fa���[��U����;6W忐�T+�оJDIֆ�?�ΒT�U��~"��ػ��Z���>�ɔ�X��?a�l�V�?Kk�#�־���+Կ�Y�|ǁ?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K[h�hhK ��h��R�(KK[��h��B�         :                 0�"]?`�1P]>�           �}@                        � �8?RB�#֭>\           �u@                        @F�&�h}�>�            `o@       	                 0��?�N��#>�             c@                        �K��?��rr��=a            @X@                        �|&�?XE(��=`             X@������������������������       �aK��H�=_            �W@������������������������       �      0�             �?������������������������       �      4;             �?
                         �Q�?S�Eo:�5>8             L@                         ����?0:�2�!>              @������������������������       �                     �?������������������������       �       �             �?                          ��?�<<0��0>6             K@������������������������       �G��'$�>              @������������������������       �O��8�1>.             G@                        �Ჯ?in�9>b            �X@                        `�?��@����=S            �T@                        ���?3q��=Q            @T@������������������������       ��Xm�d��=P             T@������������������������       �      ;             �?                        p��? ��ȓ�=              @������������������������       �                     �?������������������������       �                     �?                        �R��?�Xt�ۛ>             .@������������������������       �                     �?                        �Q�?TO�X>             ,@������������������������       ��R���>             @������������������������       �3}����=             &@       -                 P̓�?7&�%��#>a            @X@       &                 �ؐ?DF���>L             S@        #                  NA�?�F�b��>H             R@!       "                  ��M�?q��nx>=            �N@������������������������       �dX�[o><             N@������������������������       �                     �?$       %                 pM�D?F��e�>             &@������������������������       ���jF >             @������������������������       �
蕫��=              @'       *                  %+�?����0>             @(       )                 �Mn�?@�n��=              @������������������������       �                     �?������������������������       �       ;             �?+       ,                  ��d�?yZw3G>              @������������������������       �                     �?������������������������       �                     �?.       3                  ���?�H��2>             5@/       2                 Pfr�?���F>             @0       1                  H(B�?t��r߁!>              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?4       7                 ��?O�y|a�">             2@5       6                  ���?�,_��>             @������������������������       �                     �?������������������������       ���G*��=              @8       9                 �`��?-$���>             .@������������������������       ��'i�3g>             *@������������������������       �b��w��'>              @;       J                 0�/�?օ���>|             _@<       =                 p�]?E#�+��>,             F@������������������������       �                     �?>       C                 p쐺?��x��L>+            �E@?       B                 �oW�?���Ͼ�>             6@@       A                 ���?��2D��>             5@������������������������       ��lu$
U�=             4@������������������������       �      �             �?������������������������       �       ;             �?D       G                  �6�?^N��t">             5@E       F                 ��=�?�U�_��/>             @������������������������       �h�G��z	>              @������������������������       �                     �?H       I                 ܬU?�p�>             2@������������������������       �                     �?������������������������       �t��[=s�=             1@K       N                 P�!z?WE=/B>P             T@L       M                 �vu?V8���d>              @������������������������       �                     �?������������������������       �                     �?O       V                 @L7�?�Iϳ�	>N            �S@P       S                  �P��?@:-�L�=             @Q       R                ����? ��"@�=              @������������������������       �                     �?������������������������       �                     �?T       U                 �@�?@:o>� �=             @������������������������       � zML�q=              @������������������������       �                     �?W       X                 ��0�?��p-z>I            @R@������������������������       �                     �?Y       Z                 ��X�?���7x�>H             R@������������������������       �                     �?������������������������       �n�QӀ>G            �Q@�t�bh�hhK ��h��R�(KK[KK��h �B�  �:���(�>��X�C�þ}"%3�>p���5��>!ᛕ��Ⱦh ��³Ҿ�t�2࿾D�u�U�;�V�?�t�ډ��> �P&�+?�me�V�?p��5V�?�v��R��>G#<ĔU�~ڇ`��?6hA�_�׾�5wY��AO���ྊ; @�� �Ft�U�?CV�:���҈!�U�{FL�U忇�R����>��@3V�?��C#��>%�8yD�?\e6�]�Ͽ0=]j�f�ʥF�|�Ҿ0撹#h⾽	�ZԾ���J�ѿz����U�?��� �����U忚#��7Z��FJ|? �~7@!?մ#V�?r^£�U�?ߐ},Av�>�h-fU�KT
^�U�?���@���d��9����L��'啲XU�À��U忠�#�V忔��������/�[�6!�V�+GMj�U�_S?·�qĖ&@�Jy��?�vM��>Q��u��>����V�?l,.�.�>v�lkH�>­�1��>P��5�?Ϳ�ϹU�?�s,y�U忞�W�a ?��<JB�?@���U�?�� �]V�?U�N5��>��^D�U�?vvswU�?���N֑�> `�:��?����[U�?O)_?�U�?Q��P��>����xz ��
��I����x��U�\~L�U�{;��������lwU�H��T�U忦�+�1��>�k�:�U�?w������>x�)�U�?WG
���?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KMh�hhK ��h��R�(KKM��h��B�                          P��S?4%�D�'>�           �}@                        `��? T�-d�>             9@                        Э�L?C8"�;/>             7@                        h�[�>���}��=             (@������������������������       �                     �?       	                 eni?c6i����=             &@                        �4Aa?����q�=	             "@������������������������       �&=�E��=              @������������������������       �      ��             �?
                        �闾?XKO\���=              @������������������������       �                     �?������������������������       �                     �?                        �3M?`��@>             &@������������������������       �                     �?                         ����?��z��=
             $@                        �5?L�JvV~�=             @������������������������       � �-�ἅ=              @������������������������       �X�T{�=             @                         �{��?�|����=             @������������������������       ��]�=             @������������������������       �      �:             �?                        �.�?��H$'�>              @������������������������       �                     �?������������������������       �      �             �?       0                  ����?�yZ�>�           �{@       #                 ��H?�b�6{">           �p@       "                 `%�G?0@Y�%l(>�            @g@                         ���?#<r�'>�             g@                        ��??��k�.�&>�             e@������������������������       �'(J�i'>�            �b@������������������������       ���?�8>             4@        !                 P�VA?�Ɣ�,>             1@������������������������       ��� |>             .@������������������������       �p����>              @������������������������       �      R;             �?$       )                 ��,b?d��FD>S            �T@%       (                  �3��?�"�à'>             @&       '                 H��S?f�;���=              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?*       -                 .1�?%W+��=P             T@+       ,                  `��?�z5~Wa>             8@������������������������       �<>�+��>              @������������������������       ��A�����=             6@.       /                 ��?{���?��=8             L@������������������������       ���{�>             @������������������������       �n�s�=2             I@1       >                  ��?����>�            @f@2       9                 `Fe�?�*_ʗ�=             0@3       6                 X[cp?��M�>�=	             "@4       5                 `f�?S������=             @������������������������       ��GSs�=              @������������������������       �                     �?7       8                 �}�G?�X<���=             @������������������������       ��k���]�=             @������������������������       ��x����=              @:       =                 �T?P�~�=             @;       <                  0p��?@��C��=             @������������������������       � ��>��=             @������������������������       �     �׺             �?������������������������       �                     �??       F                  @��?ypQ��Y>�            @d@@       C                 p�0�?N�{�>�            �c@A       B                 p��Y?͚�wP>Z            �V@������������������������       ����s>5            �J@������������������������       �#�%y� >%            �B@D       E                 ��?��_T��=D             Q@������������������������       ����G��=             @������������������������       ��и╆�=@             P@G       J                 ���?�i)�e�>             @H       I                 ��'�?0���n��=              @������������������������       �                     �?������������������������       �                     �?K       L                  ��u�?\����M=              @������������������������       �                     �?������������������������       �                     �?�t�bh�hhK ��h��R�(KKMKK��h �Bh  D]���c���VV�w�l� �) �;��>$ճcvU�?Z �/i��>'JЖk�K>W@���?{׶�iU� ����)�>,|�,|U�?�ޮB\U�?�8��U���̛��U�ҝ>�	���W�z�~����U���uU忹q5g��Ӿ��G`U�^	}�[U�?D�5n������U�O��.U�/~��*��>�n�x���>S����>2ƥ�D��>��8I�>7����?_����ۿ?��X ?9�I�|W�?N��/V�?V��7%V�?j)�mm�վ�uumB�?H*c���>�#�#oU�?I�jU�����U�?N^K��7ܾ-{ 
��oC�N��?�j'�����R̾T.%(��?R!*ztU忖A�&��о�w��w�>�q d�{�>M��u�������\Ϳ��_3�U��]ŒTO�>c@����!�b��U�?%I˖�x�>�ꪻ��>�a lrU�?�߲^U�?����U�?���nѥ־m��+��پ5wapu��b)y��ٿ�  H��?�Hh�Ѧ�� ��U�?H+��Qݿ4BP��> �/�	?�yӪU�?b�l�U�?[̝�����w�ZUU�,؅�UU忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KKh�hhK ��h��R�(KKK��h��Bh                          �`>R??���>$>�           �}@                        `�d�?��~�>             7@                        Э�L?smX��3>             5@                        h�[�>_��n��=             (@������������������������       �                     �?       	                 eni?�o�b��=             &@                        �4Aa?��箶��=	             "@������������������������       ����b�=              @������������������������       �      ��             �?
                        (߉?6�hn$�=              @������������������������       �                     �?������������������������       �      ��             �?                        �3M?�>3���>	             "@������������������������       �                     �?                        ��?�C����=              @                         �0�?�U�p�=             @������������������������       �  <6X�z=              @������������������������       �      ��             �?                        N��S?@��ˍP�=             @������������������������       ����fዒ=             @������������������������       �      ��             �?                        ȱ�?��qà�>              @������������������������       �                     �?������������������������       �                     �?       2                 ����?Q�|�T�$>�           |@       )                 �<�?)�8�8'>5           Ps@       "                 @F�m�MS��&>/           �r@                          +Y�?$J��])>�            �c@                        ��?�^5��'>�             a@������������������������       �O��\�a&>h             Z@������������������������       ���M�>Y'>              @@        !                 �B�O?y�V�y->             7@������������������������       ���MwAf�=              @������������������������       �h4x�il0>             .@#       &                 _5?�n�&��#>�             b@$       %                 �/�?�K�M �">?            �O@������������������������       �AH\>-            �F@������������������������       ����B">             2@'       (                 P�~�?}�Ʃca#>Q            @T@������������������������       �S0J�q">             7@������������������������       �*$��}�!>:             M@*       -                 ���R?�Ÿ��>             @+       ,                 ЇW�?���%:�=              @������������������������       �                     �?������������������������       �                     �?.       /                �Yb��?"G���s�=             @������������������������       �                     �?0       1                  �ŧ?`Z
1�=             @������������������������       �  P�p��=              @������������������������       �     �к             �?3       <                 p��?3��Rg�>�            �a@4       9                 P���?�Ď	�!>             @5       6                 ��v�?��Qȹ�=             @������������������������       �                     �?7       8                 �q�?����4I�=              @������������������������       �                     �?������������������������       �     ���             �?:       ;                 ���?����=              @������������������������       �                     �?������������������������       �                     �?=       D                 �tG�?%z�'�>�            �`@>       A                 �@�?�NH���>             ,@?       @                  ?D9.p���=	             "@������������������������       �8�x�X�=             @������������������������       �$��[�z�=             @B       C                 hI�P?��>"r2>             @������������������������       �Pc�؈"�=              @������������������������       �p�ZE8��=             @E       H                  ��?�ӫG�~>y            @^@F       G                 x��?>��n�">I            @R@������������������������       �;F�� >H             R@������������������������       �      P;             �?I       J                 �%�?x�-w�>0             H@������������������������       ��Kfܲ�>             @������������������������       �D�%�  >+            �E@�t�bh�hhK ��h��R�(KKKKK��h �BX  �:�1�f�a�4����>gm�O��>ë����Ѿ��.vU�AY�u��ľ��A@��>ݶ��]�����jU�?Ղ!
���č;{U忼j� \U�r��:� ?��g�U�? 0Yv\�>���e;?D�d�U�?��{(iU�?����=f�>�i�aU�?�~��nU�? 0��j�?a��U�?%B���U�?.t8�쎬��K�~Mʾ<f�1¾�7X4�(�>����2R����P�`Լ?<����ҿ`�)o�>dK�~U�h�$�-T�?��;a�}��.V�����t^y�Ŀf�){����@�U���(r�ݿ���x���?c�Og>�/y�	ϡ��㑺�U���8� V��9#�w��H��ģU� "��\�
+�tU�rZ?VU忆 ����>��)�PE?��1��>���ҖU�?UjcV4��>��$�kU�?�9�jVU� ��C�4?|%N��U�?���5V�?�Z�����>�93]KI��a�Wwվ����1nU�?5D��oU忥��gw��:��U�]��7�U��3��+��>m��
�>��Ճ,}�?k��EV�?��6�4־L��ҳU�v��WZ���t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kch�hhK ��h��R�(KKc��h��B�         0                 pY7e?l\�	>�           �}@                        @E��?��V�9�>h           �v@                        �b'�?U�lE>(           �r@       	                 �\�?��7>W            �U@                        ���?fO�S�=K            �R@                        p�x�?�Ӫ����=J            �R@������������������������       �j�"�=F            �Q@������������������������       ��
��M>             @������������������������       �      ;             �?
                         ����?���<[-">             (@                        p���?{$:��=             @������������������������       �2C�#	��=             @������������������������       �      ��             �?                         ;��?�dr�1$>             @������������������������       �                     �?������������������������       �@16U��>             @                         ����?�z1EUs>�             j@                         ��?����=�             c@                        P�$�?��@�f��=�            �b@������������������������       ���OT�u�=�            @`@������������������������       �s�6=>             5@������������������������       �      #�             �?                        @�C�?�W��N{>9            �L@                       �R0�?6vj�B'>             @������������������������       �4ٟȟ�>              @������������������������       �                     �?                        `�ۊ?��<��>6             K@������������������������       ��0x�V>             8@������������������������       ������4>             >@       '                   .p�?�����.>@             P@       $                  �"�?��JB�>             (@        #                 x�z�?�x�z���=
             $@!       "                 �:��?E�Ȗ�=	             "@������������������������       �FO?��_�=              @������������������������       �      ��             �?������������������������       �      ��             �?%       &                 0Sf�?#��"C,>              @������������������������       �                     �?������������������������       �                     �?(       )                  @?��?2L��w%
>4             J@������������������������       �                     �?*       -                 `s5�?0�@7>3            �I@+       ,                 �$I�?nՎ\�>             6@������������������������       ���Q���=             @������������������������       �����h9>             3@.       /                  ���?���O��=             =@������������������������       ���@�1��=	             "@������������������������       �pë$h�=             4@1       F                 �2��?; �gI|>p             \@2       ;                 P n?JO,
T�=(             D@3       :                 Ў m?@�G��>             @4       7                  +i�?���=             @5       6                    �?����=              @������������������������       �                     �?������������������������       �                     �?8       9                 r'²?��vX��=             @������������������������       �                     �?������������������������       ��p��.@�=              @������������������������       �       ;             �?<       ?                 ���t?���Y�g�="             A@=       >                 @�q?�#X�8�=              @������������������������       �                     �?������������������������       �      �:             �?@       C                  ���?o}�����=              @@A       B                 ����?����\�=             2@������������������������       �                     �?������������������������       �fRnyt�=             1@D       E                 ��؈?sȭ(��=             ,@������������������������       �h1#�&��=             @������������������������       �8�y�K�=
             $@G       T                    �?1��bj>H             R@H       M                 @W�?��RO��=              @@I       L                 ��z�?�Lͤd0�=             0@J       K                  s5�?~6m�&�=             .@������������������������       �x��9�=             @������������������������       � �aqӻ=             (@������������������������       �      �:             �?N       Q                  ���?��U��=             0@O       P                   �x�?@����m�=             @������������������������       ��B4G'i�=             @������������������������       ���le��v=              @R       S                  ���?�uYN�%�=	             "@������������������������       �m�k�_=\=             @������������������������       � 9�#߷T=              @U       \                 ����?1X�w[>(             D@V       Y                 �O�?N��i��!>	             "@W       X                 p���?�h����=             @������������������������       �A.��c�=             @������������������������       ��J���и=              @Z       [                 ��ќ?���>             @������������������������       �                     �?������������������������       ��W�n�W�=              @]       `                 �:�?w��kt~>             ?@^       _                 Ш��?�x�l+�=             *@������������������������       ��j���=              @������������������������       ���� f4�=             @a       b                  �j�?��h���>             2@������������������������       ��-H�>             @������������������������       ��!q�9�=             (@�t�bh�hhK ��h��R�(KKcKK��h �B  ��ؚ;�>��5������'q�þ�>��8�>&�XXW̼��=�Ⱦ�C�� տ��=�U忄8
}�U�?��45c�>� ��r��<^�&hU�:���wU�?&|�N*?�ج|U�p����?�l�9ЪҾM���󻾑1�~������M�ӿտ��j�?7J��U�?�������|쓀��{�F�U���V忔�w3��⾇�kخ?r+�%㿜�Wx��>?W�%=�9�G��fҾ�����پ�g��^U�$-�OoU�'�K�eU�?}��#����b�ahU�#>T�V�i�=j�>jjJh�U�??WI�>����f��>���j8俣�����?��-k!����2�sU����>	�?U�EӺ��>0��N�>��am��>Z��-V��> �^E4w?��shU�?�Q
_�U�?��X�̲�>�ҥ�eU����bU�?���@�U�?�!�����>���aIc�r�ZmU�_ʒ)cU� ��~���>����Su�>��VΚU�?L̊�qU�?  FB�>����wU�?��sZU�?l7k4�> ��J��>  (-��>UUn����>�Z؇~U�?`�<eU�?=�2��U�?  Ⱥ�c�>�$�*P�>�U�[[U�?�x�bU�?9�{Eꄷ>�_�WU�?��#8[U�?��|Ҿb��mQ���n$+v�>��WpU�?+TnU忪�p����E�UIlU忍�+�U��̹�3�>Pl���>q,\U�?a�riVϥ?Xg����P\�	�iT<'aU�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KUh�hhK ��h��R�(KKU��h��B�         *                 菗Q?`#䅜U>�           �}@                        ��Ɲ?mo&�"�>a            @X@                        �x?����,
>W            �U@                        �=E?�Y{ |�>K            �R@                        �$?Z?>��P�:>@             P@                        ��IL?C�ˀ?��=             (@������������������������       ���~���=             @������������������������       �"����=              @	       
                 ��g^?��U��>4             J@������������������������       ��h��J,>             @������������������������       �α5l�w�=1            �H@                        ��G?�T�����=             &@������������������������       �                     �?                        P>-l?��5u�~�=
             $@������������������������       ���>o��=	             "@������������������������       �      �:             �?                         Yz?���У>             (@������������������������       �                     �?                        ���?��:���=             &@                        8���?
9`ќ�=              @������������������������       �W��6 ��=             @������������������������       �      �:             �?                        ����?��q�=             @������������������������       �����]�=              @������������������������       �      �:             �?       !                 �G�?����n&>
             $@                         �ZL??��"i�>             @                        ȅ !?���P�=             @                        Њ�(? om����=              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �:             �?������������������������       �     ���             �?"       )                 �vQ?���K�=             @#       &                  �P�?RG�Jh��=             @$       %                 ��O?Tr�S,i=              @������������������������       �                     �?������������������������       �      @:             �?'       (                  �G? �T�5�=             @������������������������       �                     �?������������������������       � V!���n=              @������������������������       �                     �?+       B                 `��y?k�y�>w           pw@,       ;                 ���u?h����>F            �Q@-       4                   ��?7^{�8>B            �P@.       1                 ��J�?'�3L_;
>!            �@@/       0                   �P�?�02����=             1@������������������������       �r�y*q�=             .@������������������������       ���anT��=              @2       3                 �wq?���|?>             0@������������������������       �.;�\,>             *@������������������������       �����	>             @5       8                  ���?6����!>!            �@@6       7                  y��?s;Of�8>             @������������������������       � ��$(�>              @������������������������       �������=              @9       :                   �x�?�\ >             =@������������������������       �^�}�y�=             @������������������������       ����̯>             6@<       =                 �4Π?_�-H">             @������������������������       �                     �?>       A                 �ix?Pr݄3j�=             @?       @                 �c�w? �dx�=              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �:             �?C       F                 ��>}?���
��	>1           s@D       E                 ����?���
{�=              @������������������������       �                     �?������������������������       �      �:             �?G       N                 0��q?~�ZrU�>/           �r@H       K                 @Ұ�?�w�k�	>             (@I       J                 Њ�(?��Z���>
             $@������������������������       �8������=             @������������������������       ���;�#��=             @L       M                 @b�T?�;��u>              @������������������������       �                     �?������������������������       �                     �?O       R                 �༡?DL�2>#           0r@P       Q                 �v��?�	.��>{            �^@������������������������       �qҝH��>             >@������������������������       ���{>]            @W@S       T                 �X�?����xL>�             e@������������������������       ��U���w>             &@������������������������       �b���C>�            �c@�t�bh�hhK ��h��R�(KKUKK��h �B�  Q�9B����{G@N��>�!���>s�����>R{���i�>�{ֵ��׾+ʥ֨��?�He\I⿖C^��/�>�Q��c�?�(	'��?}������ƪy�U���#��۾j��R��俨��pU�?�������IU�U�A�i���⾷�/��$�>8����ؿ�t�
qU�?&��n����f��xU���:�U�&jpF���> ����	? �F��]? �xd�?k^5a�U�?�Tʟ�U�?���U�?
"�KdU�?���m��>��DiG�>  N�(w�>�A�YU�?{�s:WU�?����;�>��lU�?Nu�fU�?,N�|U�0d��Y���af�6��O�c��ؾ7���"	�>��}�V޾���)�̿�^��U�^x����>]���Z��?<��U�?�	�n&��p���w����3V��J��.iܿ��Aq�Bܾ:<�Z� �?�q�N� ⿣�LǱ��K��V忣k�������T~�
�v�|؅U���U忤(/qU�6$�VZ)k> �Ҝi?i&���U�?.e��U�?]a�$�����	+"�of�kB���𵥜�U��sE�6�Ͽ<�l����>��;]`U��yV�U�?�Nu�
�>��T�r`�>������?Q��Ll�>X�X��žPl,Z�U忚�����t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K]h�hhK ��h��R�(KK]��h��BX         4                 �$I�?�HV�>�           �}@                        )DW?�����>�           0z@                        ��Ɲ?��|ڎ>_            �W@                        �x?�SS�>U            @U@                        �=E?Ve����>K            �R@                        �$?Z?/�Ƶ3>@             P@������������������������       �z&�����=             (@������������������������       �AxG���>4             J@	       
                 ��G?IqERS�=             &@������������������������       �                     �?������������������������       ��8 ���=
             $@                        .vz?��*�!S>
             $@������������������������       �                     �?                        ���?n�<lT�=	             "@������������������������       �F��Ħ��=             @������������������������       ��I�_�=�=             @                        ��n?��0-f>
             $@                        0�P+?Y�7����=             @                        �R�־Kl�b��=             @������������������������       �                     �?������������������������       �pR��V=             @                         �3��? ��k�Z�=              @������������������������       �                     �?������������������������       �      �:             �?                        �;�?x��)>             @������������������������       �                     �?                        p��? O�"��=             @������������������������       �@�?{W�=              @������������������������       �      �             �?       '                 5��??�fwr�>D           @t@       &                 �XZ�?��qu��>y            @^@        #                 P˦�?>ĳ��>x             ^@!       "                 ��?f[g�v>g            �Y@������������������������       ��FɀKO >S            �T@������������������������       ��	��>             4@$       %                  1��?�N���>             1@������������������������       ��
��.
>             @������������������������       �Zv
0m>             ,@������������������������       �      @�             �?(       -                 �l�?^�8��>�            `i@)       *                    �?h���V>             @������������������������       �                     �?+       ,                 @@�?X�u��i�=              @������������������������       �                     �?������������������������       �                     �?.       1                 `�>d~��Ӯ>�             i@/       0                 � �?`��OA>              @������������������������       �                     �?������������������������       �      к             �?2       3                 ��\�?�v��T>�            �h@������������������������       ��:�z�
>�            �f@������������������������       ���m���>             0@5       B                 �K��?!�/�s)>5            �J@6       ?                 �C8�?
��\��=             &@7       8                 0*��?��L�=	             "@������������������������       �                     �?9       <                 ��m�?K��0���=              @:       ;                 虯�?��o+��=             @������������������������       ��Y1��S�=             @������������������������       �                     �?=       >                   ���?�k���=             @������������������������       �                     �?������������������������       �p6��y�=              @@       A                 �-f�? ���0B�=              @������������������������       �                     �?������������������������       �      �:             �?C       N                 �vQ?�@?yj >*             E@D       I                 ��?6z���=
             $@E       F                 x}%~?t�!��=             @������������������������       �                     �?G       H                   E(�?����v�=             @������������������������       � ����=              @������������������������       � �,��L�=              @J       M                  ���?P�o��PN=             @K       L                  į�?�{���=             @������������������������       �                     �?������������������������       � �v�	�<              @������������������������       ��+ @���<              @O       V                      PI8��C�=              @@P       S                 ���?���ג��=              @Q       R                 (���?������=             @������������������������       ��:m^TI�=             @������������������������       �                     �?T       U                 ��,�?�J��h�=             @������������������������       �                     �?������������������������       ��|�梟=             @W       Z                 ���E?�p�v�=             8@X       Y                 �l�?xZ����=             @������������������������       �                     �?������������������������       � ��"Az�=             @[       \                 �H�?8��H�'�=             4@������������������������       ��.�q?��=             .@������������������������       ��u ��
>             @�t�bh�hhK ��h��R�(KK]KK��h �B�  (�Wy��|�~i��J�>äEc��оZe�)�������t�Ծ=�����M��N���?`�c0ٿ�(�����>��|��U�?�SWQ7��?��<���>u9��V�?�`�V��>z��Q�����`5�U�?y	����!"2�~߾��"�Ҿ�i �gU�H�Y�WU忬_(�����AdU�L���kU�q%�� �	�~(eU��J
�	�^v�U�wr;ؽU��J?���>�5�>��>+I1�e8�>��j���>;@��i��?߆������*Imqa�`���U�(/�kN�οJ1$�U�?��2wu֯�#�H��H���U��z�3�z���]ezU�`�+�U���N��[>�2�f��
?���V�?���I�U��lO �H���5�������&l��?��e�*ݾ�2v\�������V��ES�U�/��`�羖*��E�Ǿ�D%G��?�:�^oU念j�� ��E37��U�e
f rU�ua���Y�U�� ��U�tW����ɾw�°���� 9!i ��߂�ZU�N���Y���
�|U忹KܙU�h�q�&����;x��LyjaVU��0��VU�3ZN^UU���wn�>ӱ��Q��>����I�>)l@Y\U��a��pU�? �֓}�>C�X��U�?��ݘwU�?�׺��>ξ*× iU�6�g��U�Q{~U���k��_�>�*Zm"ȿ#���?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KYh�hhK ��h��R�(KKY��h��Bx         8                 0�"]?��rxt(�=�           �}@                        ��K�?f�����=\           �u@                         �/�?S����=�            ``@                        ��n�?}XM6���=|             _@                        �=Ű?9]�d��=q            @\@                        �Ψ?��@K'�=o            �[@������������������������       �,/����=k            �Z@������������������������       ��vS ��=             @	       
                  ��?|�U��=              @������������������������       �                     �?������������������������       �      �:             �?                        `K?��_H�>             &@                       @Oz�Z?pRS�W��=              @������������������������       �                     �?������������������������       �                     �?                         1��?�n��=��=	             "@������������������������       �                     �?������������������������       �����B��=              @                        p[R�?���H>             @                        p��?r��-�=             @                        ��?����=             @������������������������       � �<�<              @������������������������       ���z|��<              @������������������������       �      ��             �?                        ��=�?�o]�m�=              @������������������������       �                     �?������������������������       �      �             �?       )                 �Q]C?u��/�h�=�             k@       $                 P�$�?��gZ�=�            �e@       !                 ��^�?�~46U�=�            �a@                         �h��?w�x�>�=m            @[@������������������������       ��+�R��=O            �S@������������������������       �#O�Q�=             >@"       #                 `TQ�?~g�0B^�="             A@������������������������       ��s��!�=             @������������������������       �$�:��_�=             =@%       (                  �G?�?n���o>             >@&       '                 ���6?3��Kpm>             =@������������������������       �M�+Z�=             9@������������������������       �F�Ҕ&�>             @������������������������       �      �             �?*       1                 @Ws�?�8����=,             F@+       .                  ���?jBW�#�=             (@,       -                 p���?��R*M�=             @������������������������       ���h7+�=             @������������������������       �      �:             �?/       0                 X?�OSl���=             @������������������������       ��;��[�=             @������������������������       �                     �?2       5                 ��X�?�G���V�=              @@3       4                   p��?��#̈�=             <@������������������������       �~���h�=             9@������������������������       ����|7<�=             @6       7                 �-�?�.�:���=             @������������������������       ���X���=              @������������������������       �� ��m�p=              @9       <                 p�]?�\�|d�=|             _@:       ;                 eA�?��h�|>              @������������������������       �                     �?������������������������       �    ��Ѻ             �?=       J                 ��L�?��Q�u�=z            �^@>       E                 0�#�?��-,#x�=Q            @T@?       B                 pY7e?H����=M            @S@@       A                 `?��(�]?�=
             $@������������������������       �Ծ���m�=              @������������������������       �N����=              @C       D                 m�w?u��p���=C            �P@������������������������       �_����=	             "@������������������������       �a�����=:             M@F       G                 ��-�?�0�����=             @������������������������       �                     �?H       I                  ��d�?�=���T=             @������������������������       �                     �?������������������������       ��q�s[�<              @K       R                  (��?C�O;K�=)            �D@L       O                 �Ys�?�A�	��=             0@M       N                 Љ�w?J��M���=             (@������������������������       ���X��=             @������������������������       �.k(t�=	             "@P       Q                  �a�?Te����=             @������������������������       �                     �?������������������������       � �*1d��=             @S       V                 �;X?C���=             9@T       U                 �,�n?0������=             @������������������������       � `ĺ(�d=              @������������������������       ���Op�^=             @W       X                 @�d�?�{�V�=             4@������������������������       �����͈=             @������������������������       ���Ҫ�JY=             ,@�t�bh�hhK ��h��R�(KKYKK��h �B�  ҫFPߪ�>v�M���Y^�A�>�KI�>)%��V���q���'��䜥V0��!��g�T�?�m������vJ�U忼�iagU忪��~��> �AbD�?	��}�U�?����U�?"D��=��>C"e��U�?��Y�>��P.�}[�>�iէ�p�>:y�8���ǫUU�!�zUU��#�qU�? ��hy�?"9�j�U�?J�S3�U�?gz[�[���"�#�f���4�J�:��	��A�;A�����ֿ3�d}U忾*���>1K��?Tc���b��S�"�y�>�T�̽�>o_8��?eH b!�?y��U�?�<�ھ1��C��꾴A?��6Ѿ���[U忻`�dU忣W<�;��rA[suU忦F��U忋��_[�о�χ�8vǾ � $`U�^n��tL�?������d�.�uU���ZU�E׬���> �B���?�+�G�U�?_J�UU�?�Fi���>�G�<V�>���/�F�>��d!��Ⱦm�KrU�~���Aٿ7��n#��>nt���?�g�5��?�N�ڈ �)I-֌U�UU��B�>��	WU�?���hUU�?)*:貱���T�Ӿ�����0�>�sg����.�^U�?����u ������\U����zU���@.zR�>  �-I��>�96�[U�?��(_U�?ff�E���>�=2�ZU�?�e1&WU�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KYh�hhK ��h��R�(KKY��h��Bx         (                 0S�r?`�i>x�=�           �}@       !                 ���p?$_�d.>�            �o@                        �$I�?���R� >�            `o@                        ����?m��<�>�            @m@                        �?h�?�3�9�>�            �b@                        @ۣ?1
)<C�>�             b@������������������������       ��;�DG>>�            �a@������������������������       �<�����=              @	       
                  �3��?����S>             @������������������������       � �⣊=              @������������������������       ��Ӊ
*��=             @                        ��^�?<(��
��=S            �T@                        �@�?�Z�Xj�=3            �I@������������������������       ���u�W�=             :@������������������������       �Z�Z�&?>             9@                          .p�?6s�8��=              @@������������������������       ��l�Q�>             @������������������������       ��d�G��=             <@                        `��?�����=             1@                        �ㆷ?�׊gL)�=             &@                         �)�?ֽ�Uo��=	             "@������������������������       �Y*S��=             @������������������������       �����63�=             @                        ���?��O�ږ�=              @������������������������       �                     �?������������������������       �      �:             �?                        ���?���Y�թ=             @                         �_�? ��J�
R=             @������������������������       �                     �?������������������������       � tO�n�/=              @                        ����?>*C��Z=             @������������������������       �                     �?������������������������       � 5�iX*<              @"       #                @n���?�|ȦU>             @������������������������       �                     �?$       %                 `Őq?`�fkS��=             @������������������������       �                     �?&       '                  \��?��2��=              @������������������������       �                     �?������������������������       �      к             �?)       B                 ���P?)���p�=�             k@*       3                 �Y8�?kG~��>d             Y@+       2                  1��?��ÆUv>D             Q@,       /                 ���6?�.�>AO>C            �P@-       .                 `��?��R0>2             I@������������������������       �;�B=O�=             @������������������������       ��ڊc���=/            �G@0       1                 �x�=?;2����	>             1@������������������������       �`���`��=              @������������������������       �fC��Z&>             .@������������������������       �      ;             �?4       ;                 Z&�?q��qX�
>              @@5       8                  qz�?X�L���=
             $@6       7                   ��?������=             @������������������������       �����&�=             @������������������������       �     ���             �?9       :                  ���?(�%�:��=             @������������������������       �@C�'�=             @������������������������       �      �             �?<       ?                 ����?�>�E>             6@=       >                 ��s'?po�w<�=              @������������������������       �                     �?������������������������       �      �             �?@       A                  ��g�?�6qP���=             4@������������������������       �                     �?������������������������       ��#�l��=             3@C       L                 0Y?������=u            @]@D       G                  ���?��y�-^�=              @E       F                 �F}�?���>G�=              @������������������������       �                     �?������������������������       �                     �?H       K                 pj��?��wZ�§=             @I       J                 �fQ?���UQ|=             @������������������������       �                     �?������������������������       �<�H��l=             @������������������������       �      ��             �?M       R                 P\?�w)�r[�=m            @[@N       O                 ���?�?;�h��=             @������������������������       �                     �?P       Q                 �S�Y?ߌY����=             @������������������������       �                     �?������������������������       �?�d�=              @S       V                 p�,p?U@a+��=i            @Z@T       U                 ���o?N1�s�=             2@������������������������       �Q��	��=             1@������������������������       �      ��             �?W       X                 ��؈?lBP> �=W            �U@������������������������       ��c��7�=             (@������������������������       ����x �=K            �R@�t�bh�hhK ��h��R�(KKYKK��h �B�  oa�����zxz���u�pyl��A��ܵ�þ8�E�������3\g�����n^���R�ǙU�3�ؘ'?�>�lq[�U�?t����t�?^ǝ�ھ����hZ�&��ߒؿr�FW���zW��>`/�ͪK�?aXGU�ۤ��0q\��>� �����>���	�&�>)�	ɿmmªn��? ���{M?���L�U�?� �Q�U�?�g`Pzо�i�Z�?޾|�}^U忀���_U�OT�_�2�����-WU�tM�ZUU忡��_���l�T�U�-)d����D �^XU�?�^��#��*�hU��2L/zU���G轹>`�Z�A�>��C.6�>����>��~-H��>�K��Ggۿ�U��-��?��,H3���D��U�=y����?�qz�U�?5���sʾ���+��W�P�v��&cU��3WU��;��U��lt�U�Ը��hU忧�����> `��P�?n�@?�U�?i��s�U�?�'��!4Ҿ�t���U�?���~�T߿�JH�Ŀ�"v�7	��*����%�WmU忄F �zU�K�bo;w=hŏ���܀U[U�C��TXU�q!B�cU忋0�#����L~s���>a�`�U�?�0;:ⅴ>��dU�?^�T^^U��?�q����meɶ��ؾ���\eU����U忋Q:\�������\U�^�W4aU忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KWh�hhK ��h��R�(KKW��h��B                           �94W?�F>�           �}@                        ��bV?IuI��Q>[            �V@                        �U�����)�W� >Z            �V@                         e	a?u�gWy<>$             B@                        P��[?�������=             0@                         �.�?p0����=             ,@������������������������       ��+�s��=             @������������������������       ��UN��T�=
             $@	       
                  @(B�? ھM�`=              @������������������������       �                     �?������������������������       �                     �?                        T�@?�	�bp>             4@                         �Ԧ�?������>             @������������������������       � B�ivV�=             @������������������������       � �wC�=              @                        `�~?�(�e9) >             .@������������������������       �q�Yĥ��=             @������������������������       �Ŗp�Ie�=	             "@                         ����?^�	ւ�=6             K@                        �C>?q��m�=             ;@                        ?Z?4��O:��=             0@������������������������       �                     �?������������������������       ��c�h��=             .@                          �P�?BW��=             &@������������������������       �0��Ƅ�=	             "@������������������������       � ��Xx=              @                          ��?D���%�=             ;@������������������������       �                     �?                        �5W�?�A!�r2�=             :@������������������������       �{k��=             &@������������������������       ���r8�=             .@������������������������       �      N�             �?!       <                 ���f? ���>}           �w@"       -                 p>�t?�����f�=             7@#       (                 �a ?Z&W�,�=             ,@$       '                  ���?_$��=             @%       &                 0�!�?�gvC��=              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �:             �?)       *                 ��R?zN@�h��=             &@������������������������       �                     �?+       ,                 �q�4?O"ۏ^�=
             $@������������������������       ����$��=              @������������������������       � X\0Kܙ=              @.       5                    �?�ViE�=	             "@/       2                 (�e8?��p��E�=             @0       1                 �Dx?��C��Ƕ=             @������������������������       �                     �?������������������������       � �uR3 9=              @3       4                 D�"�?��,b�=              @������������������������       �                     �?������������������������       �                     �?6       9                 ��@�?T��a�=             @7       8                 �/��?�SE�=�=              @������������������������       �      ��             �?������������������������       �      ��             �?:       ;                 ��?d__�"=              @������������������������       �                     �?������������������������       �     ��9             �?=       H                 �+@?@���|1>f           `v@>       A                  h��?�7����>�            �a@?       @                 ݔ?@G �=              @������������������������       �                     �?������������������������       �      к             �?B       E                 �;�?�Co)�>�            �a@C       D                 �U��?��=��>             @������������������������       �ЕYU�B�=             @������������������������       �r�!���=             @F       G                  L��?E>�N6�
>�            �`@������������������������       �`������=             @������������������������       �\у�6
>�            ``@I       P                  E ?�����=�            �j@J       M                 �r{?��f��h>             @K       L                 x�È?{��#��=              @������������������������       �                     �?������������������������       �      �             �?N       O                    �?�gk 9�=              @������������������������       �                     �?������������������������       �                     �?Q       T                 0�2�?������=�            `j@R       S                 ��nZ?Įi�Gk�=�            `b@������������������������       ��� ݜ+>B            �P@������������������������       �v_��gZ�=Q            @T@U       V                 ��F?9���o�=@             P@������������������������       ��Z���>             .@������������������������       ���	2���=1            �H@�t�b��     h�hhK ��h��R�(KKWKK��h �B�  z��-B�>��e���>��-���>���1>�>#�&�ؾ��v����>{�6�aU�?��O2Oտ�#oω��͕U忱%��U�zF����>�|���?����U�?q��'�U�?�w
�R�>q#q�ʿ��{v*�?�Eg�ǾB[x"^V�>7f�y|Ҿke�eU�?" �dU���h5�c�>�8i.��?�=t�pU�?�mmID�ؾ��K�U�iN>AҾ�v��J,ֿ�]�ku�
�+��U�?��C����cg=��	���4�޾���!%鳾��u[���>G��oVU忰ۈ	`U�?']L�cU��%�t 㾚��zU���Ե�޾�2�`U�ઢ�kU必�3����.�l���[�HT���K{-�U�났�uU�$Q��)�����U�e�J^�U�*���۾$���c���g�dU�iW<AjU忌���O!���oC�UU�b=n_UU�j�]av�>� �r��WM"��&�޽\߷U��1��U忥��8�	���F�w�>�DCĝU�?�`���?�ty>�ž[�2�U�ڪ�	����D	 `���>k���K�> ����>?�g�#�U�?.(ץU�?b�8L���>�h~�kU�?>V*+fU���WҚ�>JS�:��>zkq1��?����]��=	�Q��þ�ݦ+>.ٿ��9����?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KIh�hhK ��h��R�(KKI��h��B�         &                 p��?�%Q��=�           �}@                        0��?B{���Z�=S           0u@                        �윳?m�_.9��=�            �e@                        �9�?4X��z�=�            @e@                        pb��?f-n��=�             e@                        в��?	_e(��=�             b@������������������������       ���rS��=�            �a@������������������������       ���Q�z��=             @	       
                 �~�?:����=             8@������������������������       ���:;���=             @������������������������       ��"r*̡=             2@������������������������       �      �:             �?                       ��;�? ܰ���f=              @������������������������       �                     �?������������������������       �      ��             �?                        �\ͥ?�`!�z�=�            �d@                         �BL??,���>             @                         ����?99貼�=             @������������������������       �                     �?                        �-�? �w�_�~=              @������������������������       �                     �?������������������������       �      к             �?                        h�b?'c{�Bl�=             @                        `I�P?��Gx&j=              @������������������������       �                     �?������������������������       �      x:             �?                         h��?V���=              @������������������������       �                     �?������������������������       �      %:             �?                        P#��?
��nȖ�=�             d@������������������������       �                     �?        #                 ���?���Tl��=�            �c@!       "                 �B��?����=p             \@������������������������       �fyuŀ�=.             G@������������������������       ��26w�=B            �P@$       %                 `Fe�?�dR��=/            �G@������������������������       �Q®����=             3@������������������������       �?�	)��=             <@'       2                 ����?�G���=�            �`@(       )                    �?��.'>	             "@������������������������       �                     �?*       1                 ����?�O�A@9�=              @+       .                 x�1e?�#��b[�=             @,       -                 ����?Ff9s��x=             @������������������������       ����ڹ2=             @������������������������       �                     �?/       0                 P���?@/��K�=              @������������������������       �                     �?������������������������       �      ��             �?������������������������       �                     �?3       :                 ���x?S������=|             _@4       9                  �x?�D}�=             (@5       8                 ���?�y��b�=             &@6       7                 pN�i?a���s��=
             $@������������������������       �<��W��=             @������������������������       �P3��D�=             @������������������������       �      �:             �?������������������������       �      ��             �?;       B                  }�?LF���=p             \@<       ?                 �CǨ?�q�x �=             9@=       >                 l#��?76P%�ٱ=             4@������������������������       ���*��=             3@������������������������       �      ��             �?@       A                 �ʁ?l��$Ve�=             @������������������������       � �Ho+V�=             @������������������������       �����߫=              @C       F                 �~�?��-t��=W            �U@D       E                  ���?��b�!�=             @������������������������       �                     �?������������������������       ��6�@��=             @G       H                 ���6?�E-MB��=S            �T@������������������������       �'��c��=!            �@@������������������������       ���~;�7�=2             I@�t�bh�hhK ��h��R�(KKIKK��h �BH  �cү�*w>\�SM��>��;g����N��ͳtH޳��[��򭧾�EX^�������	�?�C�h�Ѿٺfy���T�*Q俺MH�nU�?  ^x �>ۊ/�mU�?��oU�?)!$^K�>�S���>Uh���	?��o�U�?  �I.?j��U�?�"H��U�?��t��㰾ZhR��"Ѿ:�@\U�Ӿ��YU�  0�|a�>]��ZU�?�äUU�?eJ�A�>�|`a�U�?+q�$��>���X�>gV����?49������?zU��>a/^���?8�heU�?F)A��u�����
�1�v۬U�o�$���G�d̾?i�r�Ht>O�:VU�gA��XU�?yY�_�=��$.;hU�MdU�ˤ�1�U忓��)���z�(ta�>�wy����k_�˾��l~U�]9HB�?�8��U�?�)�D�U�?���o���f��Ҿ�8�Q���OZr��Ϳ��wjU�nq-�0��P���wU�-E�`U忳`�'yW��B�ɟcg�>� ��tU�?�ny�U�?+ި��=�����4�տHFJ����?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K;h�hhK ��h��R�(KK;��h��B�         :                  @���?Z5s��2�=�           �}@       !                  �P��?A��<�=�           p}@                          �G�?C�b���=�            �a@                        P]ڒ?�hC[J��=@             P@                        `��?I�,;��=&             C@                        ���J?��g�=             >@������������������������       �G��S=�=
             $@������������������������       ���p��v�=             4@	       
                 �DȒ?U�5��J�=              @������������������������       ��_�L� �=             @������������������������       � ��O��=             @                        0o=�?br~l^��=             :@                        P��?y%��g��=	             "@������������������������       ��]��=              @������������������������       �      �             �?                          ҏ�?�:��"�=             1@������������������������       ��I;����=             0@������������������������       �      ��             �?                        �U���!�$����=L             S@                         �\�?~�����=!            �@@                        ��Jo?"E��>             @������������������������       �ϻ�
��=              @������������������������       �L�0�D��=             @                        �e_�?.�����=             ;@������������������������       ����ٍ��=             9@������������������������       ���`��=              @                           �?E����=+            �E@                        -��?R���y�=             2@������������������������       ��<q-�=             &@������������������������       ����O�?�=             @                         ���?�i@���=             9@������������������������       ��*��\�=             0@������������������������       �4r;�S�=	             "@"       +                 v��?�<���=K           �t@#       *                 �:��?k��o�Y�=�             `@$       '                  �g<�?��4y��=            �_@%       &                 �-�|?H{��2>
             $@������������������������       ���f�A�>             @������������������������       �6W�����=             @(       )                  �H�?��j���=u            @]@������������������������       �7X��n��=F            �Q@������������������������       ��1'zc��=/            �G@������������������������       �     @C�             �?,       3                 `<��?���<m�=�            `i@-       0                  ���?�k� ��=@             P@.       /                 ���?_��$�=2             I@������������������������       ��aQ�=             5@������������������������       ��UGQ ��=             =@1       2                 �^<:?�u���=             ,@������������������������       �K6BD���=             &@������������������������       ��3-5��=             @4       7                 �,Ԗ?[U�߆�=�            `a@5       6                 ��?}�݁��=              @������������������������       �                     �?������������������������       �    �:             �?8       9                 @({�?����:��=�             a@������������������������       �͋�(S��=4             J@������������������������       �T����H�=U            @U@������������������������       �     @3�             �?�t�bh�hhK ��h��R�(KK;KK��h �B�  ܇J^���Y���t����J�ͳ�>H�F���Y.���UӾ=6w!�ľ�/�/��?8 ���ؿ��E=��0���]r���fNzU� q)at��>�k[�t��>߫�Ӌ��?�;�M�U�?�7�N�þ^�L�Ukп�Gl�uU�U3r�>H� �&�>ץ��a�>?�[�%��]�6@�U�?��rE��>�=d�L��?F��dzU�U㯫[�>�X��:ɾ���ʄӿ���bU�I�o�KS�>f;H���?v�\dU���\�"��RJ�M7˾h�J�F�Ǿ+�)�Ҽ��M�D�U�N%��D�˿S�����!K��?�K{=�տ��l_�U���NY���>��wړ�>oj�M��>؟��p�?�O2v��ÿ۶�����>�mzhU�?͎IP�U�?�u�Zе��V���m��6�d�U�F��lUU忞�CU! ��0V�8������C�?����yU�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K_h�hhK ��h��R�(KK_��h��B�         $                 �y��?𢊕�.�=�           �}@       !                 �:��?�3(��=�            `j@                         �P��?Y񊛶M�=�             j@                        `L}�?N��6��=R            �T@                          �G�?X$�d�z�=A            @P@                        �m۶?�_;�x��=!            �@@������������������������       �S�y�#�=             0@������������������������       �LS���=             1@	       
                 p��?�6
�x��=              @@������������������������       �)/Q)1g�=             :@������������������������       �)q4����=             @                        �G�?.�%VR�=             1@                       �����?%u�D��=             @������������������������       �������=             @������������������������       �4�>K�A�=              @                            �?l��@�0�=             (@������������������������       �����y�=             @������������������������       ��3��F��=             @                        PFe�?��\5�=            �_@                        ���O?}z*l��=r            �\@                        `�ۊ?S	�=A            @P@������������������������       �-��s���=8             L@������������������������       �y�����=	             "@                         ��`?#�I:ߟ�=1            �H@������������������������       �                     �?������������������������       ��h	�=0             H@                        ��=�?z
��>             *@                        ��:�?�\�ӫ�=             @������������������������       �                     �?������������������������       �p�9g��=              @                         P��?�3�x��=
             $@������������������������       ��J�O^�=              @������������������������       �\b|h|�=              @"       #                 �R��?�VF<r�>              @������������������������       �                     �?������������������������       �      �             �?%       D                 љ?�Vu�|�=           Pp@&       5                  �g<�?�[o�x�=X             V@'       .                 ���4?k���Y�=             =@(       +                  ��3�?�g�B?m�=             2@)       *                 �С?f��#���=             @������������������������       ��D�joӐ=             @������������������������       ��KC�}��=             @,       -                 ��p?.�x8��=             (@������������������������       �V��Azۭ=             @������������������������       �8P����=             @/       2                 �}]�?��(��m�=             &@0       1                 �Q�?��E�]�=              @������������������������       ���1%i��=             @������������������������       �      Ǻ             �?3       4                 lݙ|?-�w�(�=             @������������������������       �                     �?������������������������       �@��ծ=              @6       =                   �P�?�b}�j�=;            �M@7       :                 �/��?��G���=             @8       9                    �?�� Hd��=             @������������������������       ����xU"�=              @������������������������       �x��b��=              @;       <                 �N��? g��u�=             @������������������������       �                     �?������������������������       � �8Ɛ�=              @>       A                  ��M�?�����F�=4             J@?       @                 ���@?�g���=2             I@������������������������       ��5W��=#            �A@������������������������       �`*鞝.>             .@B       C                 ��Ո?�')9�a�=              @������������������������       �                     �?������������������������       �     ���             �?E       T                 ����?������=�            �e@F       M                 �ڡ3?,��\���=(             D@G       J                 @ϡ?��W�X��=             *@H       I                 ˼�?��
�W��=             @������������������������       �L(?�a&�=              @������������������������       �      �:             �?K       L                 �@h�?j�1Fq�=
             $@������������������������       ���6V���=             @������������������������       � `ќQؖ=             @N       Q                 �w��?�uvӘ�=             ;@O       P                  �_�?7=��Y2�=             @������������������������       ��v��=             @������������������������       �      Ⱥ             �?R       S                  �[??�r=#B��=             4@������������������������       ��o�)cH�=             @������������������������       ���2�#�=             1@U       X                 pa��?�Z���4�=�            �`@V       W                @tɎ?2�JtN�=              @������������������������       �                     �?������������������������       �     ���             �?Y       \                 @���?Q�E���=�            ``@Z       [                 �v@�?f�xx���=             @������������������������       �?�0�=             @������������������������       ��8�|�=              @]       ^                 �<m�?�XBu�f�=|             _@������������������������       �-��A�=$             B@������������������������       �BŠ��=X             V@�t�bh�hhK ��h��R�(KK_KK��h �B�  v]��N�U>"�:$|��>��A�b�>����sbǾ�Hk-�[>){�p-o�>�<=k}��ۻ�'�?N%*�о"oL�3��G�������Jh��Ͻ��� �b��ҚU忠�vU������׾���#��?�eƃ/俏��D|�>�w,�>�&��P��>�k���?-9E[�6�?��(_�ľ��+~U�]�C��&�����!��>U�����?���_�U�?��_�U�?�-p�o	�>�;� �U�?�'��ɿ �0楝?�"��U�?�	tpU�?�!e{қ������B;������>�W��G���U����>�Dk[U忿�r oU�?�Kg�Ӿ?I��:�?���)iU����f��>�~�� b�>�N:�kU�?��]U�a�Uj�ʾ�a`U忚�@�VU�C$��!�پXE��K��� ����-�ܶ�bnU�_�_U�1��g{���<#�U���m~U�06=Ѿ\?���Ծ,[��:j�2}���?G���&�>�Ç�U�?���uXU�lZ0]��>"����>� O����>#a% s����qU�H�`U�?�[_�z1�>�yj)Q^�?�$j]�U�?kc">\���"�2�>�-u6ß�?�qs�oU忽Mw�W�Ծb��mU�D16�ҿ=�V�H	���Nw�/���p~|y�U�ҩ1�VU��[ʹY���C:Qe�F�)��bU�saNyU� �b��>���?<��H,���t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KQh�hhK ��h��R�(KKQ��h��B�         2                 0�"]?͂F��=�           �}@                        ��K�?
rVP���=\           �u@                         �/�?�G�����=�            ``@                        pִ�?$ �X��=|             _@                        ��T�?��<LS��=y            @^@                        ����?�^.qH<�=s            �\@������������������������       ���.�=j            �Z@������������������������       �E��F�.�=	             "@	       
                   E(�?���6��=             @������������������������       �  �>`��<              @������������������������       �`�<�4�=             @                        `�|�?첻A�1�=             @������������������������       �                     �?                        0��?���Ħ�=              @������������������������       �                     �?������������������������       �                     �?                        p[R�?���O��=             @                        `���?րrkw�=             @                        �闾?X�u�<             @������������������������       �(��*�N�<             @������������������������       �     Г�             �?������������������������       �                     �?                         ��d�?p�Z=�H�=              @������������������������       �                     �?������������������������       �                     �?       '                 p��?_�#�=�             k@       "                 ��?�|���=�            @h@                        �_D�?lG�>�!�=�             f@                        ��Zy?�}�ip��=�            �e@������������������������       �QE�����=)            �D@������������������������       ��Τ�8��=�            �`@        !                 `�[�?������=              @������������������������       �                     �?������������������������       �     ���             �?#       &                 ��D�?�N�4E�=             2@$       %                 P�ײ?������=             1@������������������������       ���<�y܎=             @������������������������       ���8��-�=             ,@������������������������       �      �             �?(       +                 0��?n�@��=             7@)       *                 ��k�?�I���L�=              @������������������������       �                     �?������������������������       �      �:             �?,       /                 @�P�?VכQ]p�=             5@-       .                 �
��?DPG肦=             @������������������������       �                     �?������������������������       �0tӏ¥�=             @0       1                  �{��?.<��=             1@������������������������       ��r�v��=             &@������������������������       �T�1Kn	(=             @3       6                 p�]?��4*��=|             _@4       5                 eA�?F���y�=              @������������������������       �                     �?������������������������       �      �:             �?7       D                 p��?�J8ۊ�=z            �^@8       ?                 �u��?o}F�q�=Q            @T@9       <                 ��c�?㊠�x=�=M            @S@:       ;                  �g<�?��ջ=9            �L@������������������������       �Z�d,ޭ=             &@������������������������       �����պ=.             G@=       >                  ���?���ĺ=             4@������������������������       �                     �?������������������������       �>Y���г=             3@@       A                 �O��?n3Rq��=             @������������������������       �                     �?B       C                  'B�?�_<(�;�<             @������������������������       �                     �?������������������������       ���D]J��<              @E       J                 ����?�飌d��=)            �D@F       I                 p��?8�5(t�=             @G       H                   �0�?@��]l�d=              @������������������������       �                     �?������������������������       �      �:             �?������������������������       �      ��             �?K       N                 P�!z?Ŵf����=&             C@L       M                 0��{?���b��=             @������������������������       ��`���k=              @������������������������       �      ��             �?O       P                 ����?��	k�=#            �A@������������������������       �*f.f���=             @������������������������       ������=             >@�t�bh�hhK ��h��R�(KKQKK��h �B�  [im��>�=��G(���c�⟩>o��^!؈>H$�,��x���b��{8,;�?]�4~��;Is�*��>�	�WU�n�߇eU�?UU�����>J�_tU�?  6��n�>M�ֆYU�?��bU�?���zT�>���	��>�FX_�߽wdUU�%�VUU����bU�? `��ӵ?�2#<�U�?v���vU�?��(��D6#yǸ�������K������ZN�Y_�?r���R/׿$�i=���>Z;��{U�?�ڦ�XU�W}l�!Ծ�8�Y$�Ͼ�N��gU�s��=-�ҿm���sU����[�>  `�
�>��?eU�?��$`U�?�QN���>S~�ƾ�o��_U����hؿ�����>��,�[U�?E��VU�?�r�@$�>  �DT�>�$""}U�?K"C�UU�?�$!�%��>൹�_�>q�8���>&)Z��)�>E�N@�ɿ��\�(�?&Tè'p�,'��eU�]�S�`�?y��M�$Ծ��?�pU�UU��.w>��,�UU�?~CpmUU�?��T����'=�|M뾮��=A ھA�_U�s4o�\U�]^��zU�$v1j5�>  Ζ��>�<�XU�?�D}bU�?Dp�|�>՘�O4dۿ=[�l�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K1h�hhK ��h��R�(KK1��h��B�
         *                  @��?�il��=�           �}@                        @ۣ?��}� �=�           0}@                        0�?�?�ʆz�X�=�            �f@       	                 ��X�?
��;4�=�            �e@                        p��?P��P�M�=�            �d@                        pb��?�����=�            �d@������������������������       �	�Y����=�            `d@������������������������       �     � �             �?������������������������       �      ;             �?
                        Lpώ?J�X�W��=	             "@                         
��?ȝ|A��=             @������������������������       ��Yoҹk�=             @������������������������       ��eUx�։=             @                        ���?��
��=             @������������������������       �                     �?������������������������       �Aζ���r=              @                        �)�F?��/�BA�=             @                        �\��?P�V�1��=             @                        �U�,?`�\��Y~=              @������������������������       �                     �?������������������������       �                     �?                        �Dߝ?   #'+=              @������������������������       �                     �?������������������������       �      �:             �?                           �?��B\B�=              @������������������������       �                     �?������������������������       �      ��             �?                         E�?4�Y yq�=           �q@������������������������       �                     �?       #                 P�pv?�	��c��=           �q@       "                 p�u?�h�����=h             Z@        !                 ��\�?L�@��=g            �Y@������������������������       �t�!?	�=^            �W@������������������������       ��+�Ud�=	             "@������������������������       �                     �?$       '                 �Y8�?98���=�            �f@%       &                      �YE���=W            �U@������������������������       ��%�z�=             ?@������������������������       �c?{Z�J�=8             L@(       )                 �H�9?��(6n�=_            �W@������������������������       ��0,���=             5@������������������������       ��Z��ض=J            �R@+       0                ��#+y?����=             @,       /                  @���?�X�Q"q�=             @-       .                �}��?X�G̱�=             @������������������������       �                     �?������������������������       �a<r����<              @������������������������       �                     �?������������������������       �                     �?�t�bh�hhK ��h��R�(KK1KK��h �B�  �Z߄|Sy�f�҅���5yY�>w.��ڳ�>Û\�E�>���$��>Dڼ����?(�ɃU忽9�U�?��eK?ؾ��.G����7�]U��=5{gU忏E�]we�>�_\U�?a9=XU快*v�Cj�> @�G���>  kh:��>�'�!]U�?��7�`U�?  7[��>-j�WfU�?J���eU�?  �O�^�>��I{yU�?���+rU�?���U�����L�wU���^����ᘃ"��^t=>6���d���Կ�5C�rh�?�n�o�U�[�c��F�>�$���>5bjҹC�?]?�!%�����D��z۞��׿���сп=a@OU�>�"�}j�>�2E�X�>p�Jp[U�?c��YUU応��bU�?-��mU�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KYh�hhK ��h��R�(KKY��h��Bx         $                 ����?Ѷ0��I�=�           �}@                        �<�?���F�.�=L           �t@                        �jx?V�����=F           `t@                        ���u?�4i��=�            �j@                        ����?5։�{��=�            `j@                        @���?�'ԇ�f�=�            �`@������������������������       ���n�u��=�            ``@������������������������       �@?�BSQ�=              @	       
                 �u�?D_x���=N            �S@������������������������       �                     �?������������������������       ��hS�H�=M            @S@                        p��v?`�����=              @������������������������       �                     �?������������������������       �      �:             �?                        ��U?XGp���=q            @\@                       @O�?hz�G_��=             @                        0ꀄ?���(x3�=              @������������������������       �                     �?������������������������       �      �:             �?������������������������       �     ��:             �?                        ��*?-ݙw�Q�=n            �[@                        �5W�?��u�W�=+            �E@������������������������       �\W����=             @������������������������       �Z��@�=&             C@                        p,I�?��&O�|�=C            �P@������������������������       ���n7H=�=              @������������������������       ��U���=;            �M@                        T�4@?�f��u�=             @������������������������       �                     �?       #                 ����?�e\*��=             @       "                 �7۽?�k-��~�=             @        !                    �?����	�=             @������������������������       �                     �?������������������������       ��M�wq=              @������������������������       �    ���             �?������������������������       �      �:             �?%       @                    �?�8��A�=�            �a@&       3                 Ь9�?.�����=;            �M@'       .                  �!�?U��?��=             0@(       +                 ����?����a��=             *@)       *                 ����?���5��=              @������������������������       �                     �?������������������������       �                     �?,       -                 '�,l?��K�t�=             &@������������������������       ���x/�q�=             @������������������������       �5J�\�*�=             @/       0                 ����?� ���?�=             @������������������������       �                     �?1       2                 (�?2�+��]�=              @������������������������       �                     �?������������������������       �      ��             �?4       ;                 ��[?*��z�I�=+            �E@5       8                   p��?P������=             3@6       7                  `���?�k�~���=             *@������������������������       ���<�=             @������������������������       �d\��XU�=             @9       :                  z�?�"a��"�=             @������������������������       ��3���'Y=              @������������������������       ��F��&I=             @<       =                 �࡬?7�o�M�i=             8@������������������������       �                     �?>       ?                 ��ח?�)&�QY=             7@������������������������       �x�e��R=              @������������������������       ����TG=             .@A       P                   ��?�Yg1�B�=Q            @T@B       I                 @�-�?�U�����=3            �I@C       F                   s��?� �ԫ.�=!            �@@D       E                 P��?����H�=             ,@������������������������       �菕j�=             @������������������������       �w��ݡ=	             "@G       H                 Q�?yӓ��=             3@������������������������       �+�y?��=             2@������������������������       �      �:             �?J       M                  �K�?��DCs�=             2@K       L                 ��?�B8=��=              @������������������������       �PN�K�g�=             @������������������������       ��,��{=             @N       O                 0�6�?������=
             $@������������������������       �$yi��=�=             @������������������������       �*��BZ�W=             @Q       T                 0�Ь?R�>��U�=             >@R       S                 `���? �8���<              @������������������������       �                     �?������������������������       �      ��             �?U       V                 0���?|!ʋѨ=             <@������������������������       �                     �?W       X                 @��?�d�VH�=             ;@������������������������       ��~/BS(�=             @������������������������       �^�h���z=             7@�t�bh�hhK ��h��R�(KKYKK��h �B�  v���%h�t��S�-��*�1����L�Ϙ���>
���"��>l�*������񞥿����jU忢�)���>Dd��U�?�i{	��? ��-���>�W��U�?�Ѝ�nU�?Ow�3¾�%'	t��Y"�b�����'jU��D/ppU�F�YWU快��Pܭ���z��Ѿ������?&��v��ɚ��j�����9�oU�H�[=v�?uvE��\��{�U���1O\���L����־4�[�&�޾%�܈bU�
�>^U��0�gUU忓���qU�`s�Wd��>��`l{B���C��Ҿ�y���|��  �ń�>����VU�?�2b`U�?Z_�cb�Ǿ����C�9�o�o׿�.�֣_�R[���U�/�0��bվ��v�`U必��4XU�?���ݥ>��P6�>F���C��>�(f�3�?��ƳeU�?�,�ƾ_���_U忎��VU必�c�oӨ����ZU�	�ꁤ����EWU�M�R�VU����v���>�'�L� �>��g�(!�>uWY���>�E5MfU�?{@�TKY�?}�c�T���=����¿m�O�hU�?�[�`��>���+�6�>V8_^U�?6�RTZU忮`�L$�>��6hxU�?��WU���[�9x�� �A����>B��`U�?(ڦ�`U�?���~����dU�?�C�:����o�cU�9y�XU忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KMh�hhK ��h��R�(KKM��h��B�         *                 0���?p�3��ն=�           �}@                        �6Sz?' C���=R            u@                        �r�w?��)o�=,           �r@                        ��h�?z3p!*9�=)           �r@                        @@�?�e��g�=�            �l@                        ��=�?�3�CM�=�             k@������������������������       ���7vX�=�            �j@������������������������       ���3K"��=              @	       
                    �?�k����=             ,@������������������������       �������=
             $@������������������������       �eS�+f7�=             @                         `jS�?Ih"婕�=C            �P@                         ����?G��i���=@             P@������������������������       ������(�=/            �G@������������������������       �z ڭ���=             1@                         ����?��+���=             @������������������������       ��8�j�6p=              @������������������������       �      p:             �?                        �/��?|��0j�=             @                        �ny?�_� >9F=              @������������������������       �                     �?������������������������       �      P:             �?������������������������       �                     �?       '                 P!d�?"����=&             C@                           ��?�W�G��=$             B@                        ��Q�?��P��=              @                        ԏ)�?�)�)��=             @������������������������       ��ͣ�niK=              @������������������������       � ���l�G=              @                        �ơ?\�LY�Z=             @������������������������       �                     �?������������������������       ����A=             @!       $                 ����?��9���=             <@"       #                 8,�?��[*P�v=             7@������������������������       �ؒ	�d=             &@������������������������       �t���@Nv=             (@%       &                  &&�?��%`�֫=             @������������������������       �                     �?������������������������       ������`=             @(       )                 ��H�?M�/v�=              @������������������������       �                     �?������������������������       �                     �?+       .                 @K�?�1s}�=�            �`@,       -                   ��? ��B6��=              @������������������������       �                     �?������������������������       �      ��             �?/       >                 �Q�?҆�(\�=�            �`@0       7                 �ز�?y��?#�=`             X@1       4                 �U��>�P8���=             7@2       3                 W�?�%exzf�=
             $@������������������������       �Rx&,"�=             @������������������������       ��(f���=             @5       6                  ���?0#�J��=             *@������������������������       �ſ����a=             (@������������������������       �                     �?8       ;                 p���?Q�9�ۯ=I            @R@9       :                 @��?�od/�=             1@������������������������       � �L�!�<              @������������������������       �d��=             .@<       =                 `Fe�?˪��JU�=8             L@������������������������       �<9�E��=              @������������������������       �a1dA�=0             H@?       F                 �s�?�!��ۮ=$             B@@       C                 �I�?hXnS�a�=             8@A       B                 v�؁?�;G� r�=             6@������������������������       �K��4D�=             2@������������������������       �`�#���y=             @D       E                  `�J�?�T�(�d�=              @������������������������       �                     �?������������������������       �     �b�             �?G       J                  ��^�?��]�dj=             (@H       I                 pX��?,��S|i=             @������������������������       �(@G�ь2=              @������������������������       �В1QӷW=             @K       L                  Ή�?>���Jh'=             @������������������������       ���ڒ�=             @������������������������       ���'�
�<             @�t�bh�hhK ��h��R�(KKMKK��h �Bh  �Bg���>�+��w��Hg�F�󕾆=�������V�&�M��cQƒ\����wO�Iֿg�օy(�?=�5��v�>�Eҗ���?W�K��2�?�4̆�ѳ��(E���s����Ŀ�U�3��߿o>���>�vfU�?���ZU忯�=�־@tB�~6ƾ��O�YU�%��zXU�b��dU�d@��.�> ��D<�>  �T	�> �P���>th�[U�?	/`U�?  ��ĵ>��3pXU�?2(�VU�?o�7ޓڳ>No��ӕ�>9���WU�?d�'<YU�?VF5��k���)�p`U�wP�JWU�?&(V�qվVlUU�?��ɷcU快9Nȅܫ> �6%�/�>�Q(+kU�?ygy�rU�?g�<�/��>+�@���>6��/_�>�Kz���>҇knU�?� �)�?�\�����>t>�� +�?��H?_U�?aބ,�>�#��:��>T|n{_U�?@�c���?I6���Q�Cv�Y��޿1�5���?��d��������¾�v�i׽���-��\U�5]��XU�?)r܎�⾺j3?nU忀�%7VU�?UU��:��>  ��6�>L5�qVU�?�з�XU�?%Iv�2�>S}x�UU�?/m�oUU�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KMh�hhK ��h��R�(KKM��h��B�                          �߯�>֐��-�=�           �}@                        �m۶?�LSV�=             5@                        �--�?vQυ���=             2@                         `S��?� 夷�=             ,@������������������������       �                     �?       	                 �jA?����6P�=             *@                         �Ԧ�?f�޽L��=
             $@������������������������       �Z��)xƠ=             @������������������������       ���5�s�=             @
                         �я�?����c=             @������������������������       �                     �?������������������������       ���p�N�F=              @                        0~��?9'����=             @������������������������       �                     �?                        P�,�?N7Ч!=             @                        ʊ�X?i̌ ?=              @������������������������       �                     �?������������������������       �     @�9             �?������������������������       �                     �?                           �?��7,*�>             @������������������������       �                     �?                       ���Ou?��<�:�=              @������������������������       �                     �?������������������������       �      p�             �?       2                 p^�e?}���@	�=�           0|@       #                 0�G?H�6���=0             H@       "                 0��m?$*}���=             6@                        �<��>�/'�E��=             5@                        �)�*?�S�c���=             @������������������������       �                     �?������������������������       �  �Ӯm�<              @        !                 `�]?y�F���=             2@������������������������       �gɐ�L�=             @������������������������       ���ha�=             &@������������������������       �      Ⱥ             �?$       +                 ���`?��^9߭�=             :@%       (                   �G�?�F��t�=             0@&       '                 p�1�?`f�=             @������������������������       ���=���=             @������������������������       �     ���             �?)       *                  �~��?�3���=             &@������������������������       ��s��8��=             @������������������������       ��$w�R�=             @,       /                 `��?T��I>(�=
             $@-       .                 ��qb?�x�����=             @������������������������       �                     �?������������������������       ��\����=             @0       1                 ���@?�"��=             @������������������������       �Ф7���=             @������������������������       ��ɒ8ٕ=              @3       >                 ��l?[gV9_�=�           0y@4       7                 #~&?(�'&�=	             "@5       6                 ���i? �5�&V[=              @������������������������       �                     �?������������������������       �                     �?8       ;                 A�n?R�Q�=             @9       :                 �+�k?<�eT��=             @������������������������       ��.��e�=             @������������������������       �                     �?<       =                 ��dt? �9P.i=             @������������������������       �                     �?������������������������       � �m`�?5=              @?       F                 0'Fx?�c��@N�=�           �x@@       C                 ���u?۰�O�=%            �B@A       B                 ���>J1�꛺=             ;@������������������������       �                     �?������������������������       �+�*�>�=             :@D       E                 ��G�?�(��3�=
             $@������������������������       �X�,@���=	             "@������������������������       �      �:             �?G       J                 �To�?]����=e           Pv@H       I                  �Ԧ�?���%�=             >@������������������������       �                     �?������������������������       �F�~�K�=             =@K       L                 �m۶?���c��=G           pt@������������������������       ��Q�;梾=5            �J@������������������������       ��1y�X�=            q@�t�bh�hhK ��h��R�(KKMKK��h �Bh  >����_���tQ��ɾ�{��e��Ӧ�?x2�>����`U����ټ>
����M�>X��7^U�?e�Yw���?sq��@���X�� VU����XU忢�*�Uݾ��Q�{U忨��B�����1*�}�Y���UU忇�rZUU忮R��UU�]�ǟX��ܠ��U�r9����>IC�[U�?�z��ZU忘c�i�}>���}��>���Pݰ�@�V��k��4�.۾���ZU忓���`U�zWD;c�>d�����?��d�ӿ�=\nU�y� �8��>0XN���>b�6�(�>O.M=eU�?�i-�UU�e���sȾҠwbU����B67�?�n	���>�hJ�޻>�5}]U�?�,�6&�?�*n��;�>I�gU�?��tU�? �N��y�|a�7�b�������Z��@pU��&��qU念'-�!tԾ�G�zN����p2�X����*_�\U忯��1������7dU忏S�aU忕�)��w>�q�Y��>�"1Nq&�>JRUgU�?8���	�s�Ӥ޵��>�����?Aey�xU�?�es�o,���X�"þz.%sU忌m���Ϳ�"J��~p>R�S���ؿ@e��JѴ?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KKh�hhK ��h��R�(KKK��h��Bh         *                 �94W?;EF�c�=�           �}@                        �U���d�����=[            �V@                         e	a?�GE_��=$             B@       	                 �$?Z?g��|��=             0@                        pF�T?��
C�=             *@                        ��N?Hpi$�ծ=             (@������������������������       �f3�ƏP�=             @������������������������       �P�O(�ß=             @������������������������       �      �:             �?
                        �Q�?@\`oT0�=             @                        �؉�?`I���=              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �:             �?                         �%c?���p�=             4@                         �JV�?��f��\�=              @������������������������       �                     �?������������������������       �                     �?                        �aH�>.�_�(��=             2@                           �?�O/���=              @������������������������       �                     �?������������������������       �      ��             �?                         ;��?��,���=             0@������������������������       ��b�igg�=             @������������������������       �u�El5��=
             $@       )                 ��bV?���I��=7            �K@       "                 P^N<?ՙ���ٳ=6             K@                        `��?-l��=#            �A@                        `�լ?�w��9�=             0@������������������������       �pf�k=             *@������������������������       ����L7X�=             @        !                 ��-?ONݥŭ=             3@������������������������       �rڎ1ш=	             "@������������������������       ����=
             $@#       &                 ��V�?r��P�ж=             3@$       %                 ��j�?�DlgD�=	             "@������������������������       ���qZܣ=             @������������������������       �{w6�1�=              @'       (                  @(B�?��1�$�=
             $@������������������������       ���5��p =             @������������������������       ��#Ҷ�w�=             @������������������������       �      �:             �?+       8                 ���h?�����=}           �w@,       7                 �M�h?bV��q�=             =@-       2                  �\�?d_-���=             <@.       1                 `��?�����=             @/       0                 @F�@,TV'�=             @������������������������       � s3�e�a=             @������������������������       ��,�m]�b=              @������������������������       �     貺             �?3       4                 P+�Q?(��1�=             6@������������������������       �                     �?5       6                  ;��?��s�s�=             5@������������������������       �0<{֥w�=             0@������������������������       ��f�7��}=             @������������������������       �      Ⱥ             �?9       <                  ��i?�$��8�=`            v@:       ;                 �U�,?X���=              @������������������������       �                     �?������������������������       �      �:             �?=       D                 �To�?h� �=^           �u@>       A                  ���?���Ϙ��=;            �M@?       @                 0���?�����W�=)            �D@������������������������       �ٛ|��3�=%            �B@������������������������       � B˞)�=             @B       C                 ���H?�#-FJ��=             2@������������������������       �������=              @������������������������       � ?"Jm,�=
             $@E       H                 ��n�?ad�7Q�=#           0r@F       G                 z�?�4_��=�             `@������������������������       �MCzI���=             9@������������������������       �Ś����=h             Z@I       J                 ���?�(nz���=�            @d@������������������������       ����e}��=             (@������������������������       �`�{/�=�            �b@�t�bh�hhK ��h��R�(KKKKK��h �BX  �L8\��w��Z����>߇�1�&�>��hW����i�c%9�>�Ru6�;�>��
��?��^U�?���{bU�_)�]���R�f�辉��hU�4��bU�{'�xU忾���Z��> ���l?⅐~nU�?���4�U�?R�T�/n�>�Sl�cs��^�\U�vM?�eU�_=�rg|�>)%��pU�?Mr���s�?N�ĭ��Q)��͵�tC��ƾE��n���5zXU�_k��@�?Jw�G٢о��"ZU��9BZaU�ur��V�>$=@'��>Qoe�_U�?Z��F�<��i!,����/��VU�?�o�[U��� =sU�?QrVV�>���SV5�о���W;T����\@]�Q�V?eU忮,6@aU��lVU�H)�ٟ��,�"z]U�?�7�Z�ľ�"i�xZ�^�u��?/ݡpU��Br�ux��Y�����>[��6~U�?o��WU�,�������ǋp��a�>񜔋�V�>z���?�P�gjU�?I�Dt��X4ڡ w�2"�	���?v�H���=
cp���#����;ۿ��V�����/t�Q��>S5���?��Τv��t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kch�hhK ��h��R�(KKc��h��B�         (                 �r��?0�����=�           �}@                        ���?2�%d��=�            �b@                        ��6�?�X��=�            �`@                        ��5�?@_5���z=~            �_@                        P^��?���.)�n=y            @^@                        �zۦ?ء��pS=q            @\@������������������������       �"���0O=p             \@������������������������       �                     �?	       
                 @F�E�;ea�=              @������������������������       ������h=              @������������������������       ������=             @                        �'��?��J��=             @������������������������       �                     �?                        �b'�?� �{��=             @������������������������       �x���&�O=             @������������������������       �      `�             �?                        H1�r?j��M��=             @                         P�J�? �-�c�B=              @������������������������       �                     �?������������������������       �      �:             �?                        PJ�?Jp����r=             @������������������������       �                     �?                         �g<�?T�v�W�P=             @������������������������       �                     �?������������������������       � T����<              @                        �7?E�7ƙ=             2@������������������������       �                     �?       !                 p�:?��͸��=             1@                         `���?/�ܥLR�=             &@                         `��?���Ȫ��=
             $@������������������������       ��A�y�4Y=              @������������������������       �4���$��=              @������������������������       �      ��             �?"       %                 @W�?d��x�Q=             @#       $                8��t�?��#N^2=              @������������������������       �                     �?������������������������       �                     �?&       '                 �m�?�*�+*=             @������������������������       � �IG��<              @������������������������       � m<:�Ơ<              @)       F                 p�v�?�
���=B            t@*       7                  ����&����=v            �]@+       0                 0{��?;%;���=&             C@,       /                 �y�?!E��%�=             0@-       .                 �J�?��R�L(X=             .@������������������������       �<��ڷx=             (@������������������������       �| >q|�d=             @������������������������       �      ��             �?1       4                 ��Dm?��7A��=             6@2       3                  �d%�? �0߃��=             0@������������������������       ���͞��=             (@������������������������       �Yi�~�u=             @5       6                   \��?�X�z�=             @������������������������       ���lXp��<              @������������������������       �@0e?juz=             @8       ?                 �<�?���B]�=P             T@9       <                 �\��?*Z�cl�=              @@:       ;                 ��p?7)���ƀ=             >@������������������������       ��X���Qy=             5@������������������������       ���&��}=	             "@=       >                 hs5�? ���F=              @������������������������       �                     �?������������������������       �                     �?@       C                 pM�D?(7�w�=0             H@A       B                  �P��?eV���=             @������������������������       ���H,B�{=              @������������������������       �                     �?D       E                 ���?
�ʉ��=-            �F@������������������������       �                     �?������������������������       �,Z���i�=,             F@G       V                 ��|�?*��a�S�=�            �i@H       O                 Ц��?Z���4x�=^            �W@I       L                 ��?��]�}�=A            @P@J       K                 ��`�?j^/��e=,             F@������������������������       �4�����M=!            �@@������������������������       �;C�ޱ1w=             &@M       N                 �p�?� +l�E�=             5@������������������������       �^i���S�=              @������������������������       ��L8$)�=             3@P       S                   .p�?t;q�=             =@Q       R                  ��?QjQnK*�=             @������������������������       �BXh�\,B=             @������������������������       �      �:             �?T       U                  @?��?b�O�`�=             9@������������������������       �                     �?������������������������       �yv�H�v=             8@W       ^                 `WJ�?�@��,�=n            �[@X       [                 г��?�3"d���=             3@Y       Z                 ��>�?x��2�t=             0@������������������������       ��<|��	j=             *@������������������������       �NA87�Pq=             @\       ]                 ��x�?�Ыӛ�=             @������������������������       �[�+�-|=              @������������������������       �                     �?_       b                 @8��?�t\���=[            �V@`       a                 �5Ry?�c ���=Z            �V@������������������������       ��S�ꠔ=1            �H@������������������������       �┑��օ=)            �D@������������������������       �      ��             �?�t�bh�hhK ��h��R�(KKcKK��h �B  �O��c�>q�),#��t��]R���մ���b���tl�:���P�_F���� �VU���1�XU�? ��c���@_�\U�<��U��^g���>���`U�?S�C��눾�!�WWU�FR��YU�?�Q�T���>  �C�>|���]U�?�7!�^U�?�+T�4��� �IWU�?+8*�������|UU忤"�VU���{�eϸ�ɍK�aU��D�h������^�3��*G�'�1�����WU忐hn}[U忿��\U�u<���[|>T��k�����Qx�UU��UmVU�   ��O�>t�9VU�?x�̟UU�?��mA��>��j˖�>�COoo!�>��bp�n�޿�A8՜�kG�UU����WU忋=]U�?n"e-��>D�ִF��>�W
��?�"x�+8�?G���&ž���UU�t��[U�μ��;�>���]6?��,A����p�1̈́*�?��n���y�1�JӾ��RS\U��3[U���;[�Ұ>�~œX��>��E���?Z��iU�?�D�b�(�>��W_U�?GB�>��?���Q�z����at���wḶE竾�8�\���w��ߏܿ�� �t��]	n5��'&�ecU�%�.Z}s߿Ȩ���]�>*ޛ��2;��.qVU��t�nfU�H#o9��>ͱ%�_U�?�}�c`
�?!K����>��/����>���i�>?tc�/�̿���PXU�?���m�I�>q����?o�,qU�?r},����~��&�s��Hѿ��2g���?�>�\^U�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KUh�hhK ��h��R�(KKU��h��B�         *                  ���?y#�rB��=�           �}@                         (V�?���C�=4           @s@                        ��{�?<m����=,           �r@       	                 @�?�7�	��=f            �Y@                        ���?nP����=4             J@                        �e]�?�q�$�y�=3            �I@������������������������       �	�Mϡ�='            �C@������������������������       ����8�_�=             (@������������������������       �                     �?
                         ���?,}�ę/�=2             I@                          ���?VQMo\֢=(             D@������������������������       �� e�ߎ=#            �A@������������������������       �
G(j��=             @                        LR��?Ʌ�z�u�=
             $@������������������������       �����s�j=             @������������������������       �C7�i�od=             @                        �&�?l,�i�=�            �h@                        pB�?N�æL��=�             `@                        �2*�?�+�!�=}            @_@������������������������       �]O���ۼ=             >@������������������������       �N�3�m�=_            �W@                        Њ�H?I�̲�x�=             @������������������������       ��D��2��=             @������������������������       �      ��             �?                        ��6�?<A<�b��=E            @Q@                        �2OF?��h�	ޜ=             8@������������������������       �"�\9��=             &@������������������������       ��t�`w=             *@                        p���?�CƝ��=-            �F@������������������������       ��ȩ+��=             @������������������������       ���5ى�=)            �D@        !                  ]`�?-'��8�=              @������������������������       �                     �?"       )                 (I��?�����=             @#       &                 �D��:I~찁u=             @$       %                 mG�?D���{=              @������������������������       �                     �?������������������������       �      P�             �?'       (                 �g'�?��vS�1=             @������������������������       ����f<             @������������������������       �      :             �?������������������������       �                     �?+       <                 0��?+�uc1�=�            �d@,       -                 0��?މwpݕ=>             O@������������������������       �                     �?.       5                 �@�?�Y�P�I�==            �N@/       2                 �$I�?|��j��=             8@0       1                 `f�?�l��=             &@������������������������       ��8|Ć=             @������������������������       � K��{�=             @3       4                 ࡭6?31kA�=             *@������������������������       ���awt$s=	             "@������������������������       � ��/F��=             @6       9                 ���?�b�9z=%            �B@7       8                 ��N�?YN�&D�i=#            �A@������������������������       �(�CT��=
             $@������������������������       �-.�j%6�<             9@:       ;                 �b'�?DaA�/�=              @������������������������       �                     �?������������������������       �                     �?=       H                 �.��?䪅sM�=f            �Y@>       E                 �2)�?!����z�=             0@?       B                 ���?!";iI�=             ,@@       A                 �G��?ܣ#���=
             $@������������������������       ���y�=              @������������������������       ���Glœ=              @C       D                 {�?�2^�/��=             @������������������������       �                     �?������������������������       ��z��]J�=             @F       G                 �+�?06UP�z�=              @������������������������       �                     �?������������������������       �      �:             �?I       N                 ���?k��Ͳ�=V            �U@J       M                 p�v�?�87���=             @K       L                  ����?G.�'q�=             @������������������������       ��@f�:�<             @������������������������       �      ��             �?������������������������       �                     �?O       R                 ��q�?���zv�=Q            @T@P       Q                 ��K�?��{�7n�=             @������������������������       �                     �?������������������������       ��.�	��Q=              @S       T                 0{��?�P�Q5�=N            �S@������������������������       � ��@�c=              @������������������������       �\��uV��=L             S@�t�bh�hhK ��h��R�(KKUKK��h �B�  �a�~3��y4��iڈ>�,B��>�
2��Q���Y?�>C�֙� �>���Q<�?�V��nԿ��gU�?�-�3 N����:�{���W*wٿ��cU忊�q����>�{ �XU�?�{}�WU��_V�â>o% ��c�>���ڰ��>|�uj���?DoN�<�?:D���>�7-�dU�?��6�VU��"��Y���"�<�¾���Q]U忸jP�XU�)�u`�>lW�P�?�U�?�b��z�þ�7cU忥��a��ٳ1�qd��x^Dm�����:<�YU忽��:VU�7�"�
��u3�WUU�k`�%VU忻S �[U忔��j�%��D��Ezv>E�f\U���1��>���I*x�>Gv���T��q���?���[U��q�>K��>���.��?�YNa]U�?�#ȋ�U��R�h�����m�TZYU���i�UU忉	jL�"Ⱦ���UUU��7t`]U���'zv��șD@�sѾ�����t��
���b>����?~M��[U�%�I�cؾ0�~�mU忝M)uF\�D�0!��������U�P��"eU���i��0��z��*�̾���o$���[���UU応%��_U忣��GbU�p���뛜�����>�X�UU��J��[U�?�lV嫁��@UJ\U�av��ѿ�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kih�hhK ��h��R�(KKi��h��B�         2                  ���?}u�K�|�=�           �}@                          �G�?�(����=4           @s@                        �7~�?��g{�=@             P@                        0���?���t�=?            �O@                        hO�?�V㿧�=6             K@                        �M}C?T���b��=1            �H@������������������������       �Fp�_Ց�=             ?@������������������������       �x�/����=             2@	       
                  �Ԧ�?_��Rm�=             @������������������������       ��,%Vx�a=              @������������������������       ���m���U=             @                        @��?�yG��,�=	             "@                        �C8�?$�_�jt�=             @������������������������       �@��u�;n=             @������������������������       �                     �?                        ���R?�M˴,��=             @������������������������       �                     �?������������������������       �B��bj=              @������������������������       �      ��             �?       #                 ��C?�����=�            �n@                        0�q�?mQN�T�=�             e@                         �P��?���^�d�=�            �a@                        �U���Ԙ�i�ĳ=0             H@������������������������       ��蕭0|�=             :@������������������������       �1u����=             6@                        @�V�?��z��=]            @W@������������������������       ��"���g�=\             W@������������������������       �      �             �?                         p�F�?�H����=             ;@                        pi��?h�}��=             @������������������������       �8-	��"�=             @������������������������       �                     �?!       "                  ���?�K��ޝ�=             5@������������������������       ���:H�=             2@������������������������       ������Џ=             @$       +                 ��K?�P.S�=L             S@%       (                 ���v?�-�t���=             @&       '                 ��sn?��Q��ϖ=             @������������������������       �Z6S�js=             @������������������������       �      `�             �?)       *                �����? ;;ȡ=              @������������������������       �                     �?������������������������       �      �:             �?,       /                  �g<�?Wn*T�l�=F            �Q@-       .                 `��r?�j��"l�=             <@������������������������       ��Sō�=             1@������������������������       ��e��l�g=             &@0       1                  X1c?�Q�Czf�=*             E@������������������������       ��Q�r�=	             "@������������������������       ����|˫�=!            �@@3       R                  ��?]�:(��=�            �d@4       C                 �T�x?�v��.��=o            �[@5       <                 �m��?w�R23�=R            �T@6       9                 ���x?����U�=4             J@7       8                 p��k?Bmy���=             1@������������������������       �xQL@X1�=             (@������������������������       ����"��R=             @:       ;                  `S��?�k;�Ȥ=#            �A@������������������������       �R4M��0�=             .@������������������������       �f��Kl�=             4@=       @                 B��?c������=             >@>       ?                   +Y�?̼�q�=             1@������������������������       �x����=
             $@������������������������       �]Z<�s5�=             @A       B                 ����?ڠz�>�=             *@������������������������       �����Ě~=             @������������������������       ���hK�t=
             $@D       K                 p'�?X�rBD�=             =@E       H                  �_�?���|X�=             6@F       G                 �A��?�5-F�t=             *@������������������������       �@�Uj#K�=              @������������������������       ��~��)B=             &@I       J                  `<��?V�>�	�=	             "@������������������������       � ���%:=              @������������������������       �P�ss=             @L       O                 Pc��?�{P�&��=             @M       N                 ����?0��<�g=             @������������������������       �                     �?������������������������       ��ƶ1E|M=             @P       Q                 �sW�?:��j��b=             @������������������������       �                     �?������������������������       ���ȌG=              @S       Z                 ����?�=��'�=5            �J@T       U                 Pe �?8FK+���=             @������������������������       �                     �?V       Y                 Pez?i��6j�=             @W       X                 ��i?��ȣ�=             @������������������������       ���`�<              @������������������������       �                     �?������������������������       �                     �?[       b                  (��?#��4�=0             H@\       _                  �E�?�M� �=             =@]       ^                 �j:�?㑪lu`�=             @������������������������       ������=              @������������������������       �k��u���=             @`       a                 @4��?Z<���=             8@������������������������       �ZT�L��=             1@������������������������       ��~�K:�=             @c       f                 hx�_?��_��z=             3@d       e                 @|��?�����=              @������������������������       �                     �?������������������������       �     �H:             �?g       h                 0o�y?D��=��3=             1@������������������������       ��0^ޮ=              @������������������������       ��w��.w=             .@�t�bh�hhK ��h��R�(KKiKK��h �BH  �T��P5u>ڑ^ϪF�����v���>�ILϣ>y� 4���>�]��>V߱��?C�+4���$�z��ʾ�	d^U�O��\WU�=�4���>  ���p�>�`�`ZU�?Z��`U�?�{�?[F�>=�FXU�?P)4�WU�� �1cU�?w')i~͞��bʢz���	ӷ������k���R��߿� \o)������՛>�:sE��?Ac�fU�?�|E��Ⱦ9}��d徺N?�aU����wU�c�P�7e��޽ Z}��D��]U忢 �����>���_�%�>їb(h��>IH��XU�?ߤi�YU� �\E��>jJ��oU�?=)hU�?[�w� 0��k�+�ƻ�>l��YU�?�<�F��ҿ�e䩄f��+o�࿸h��{�����2��>}��|Z~>r��J��>�l:q����FD���>52��u2��+v��[U�?��q��x���Z<O㿲��=���?D	G*��>�8��O��>V�B|�^�?@50�w�?���zo���n��ZU�C�5����?@��#�g��9iq���Y��
	����߸ZU�k(ZVU�t���9|Ⱦ��]U���XU�5���&D�>  �`��>!iq�YU�?{�Z�WU�?0Z�H��$��WU忘�O�UU�6�� _�>�Z�V%�>�0�U�?ώ�@:��>s49�~��T	�gUU�w��UU忺���eU�?��u$���>���h��>��a$��>EA�fU�?]��i�V�?E��TU��>��]�y����4����?�V��$���p&��Ǿs�/]U��*zUU忏�`�L���%G�VU�2��UU忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KUh�hhK ��h��R�(KKU��h��B�         &                   s��?�y�#҈=�           �}@                        pҷ?�)ݷ�w=�            �e@                        ��e�?���h=w            �]@                        ��ё?��c�$[=o            �[@                        (/��?��7�U=k            �Z@                        p(�?j�G�B�P=i            @Z@������������������������       �@L��	I=b            �X@������������������������       ���Ta=             @	       
                 �'U�?��Ku%�=              @������������������������       �                     �?������������������������       �                     �?                         ��3�?��O�3p=             @������������������������       �                     �?                          ��?��l�;=             @������������������������       �                     �?������������������������       �=�⛘ =              @                        ��A�?��|�=              @������������������������       �                     �?                        0vb�?sH2�q>n=             @                        �j��?���^�8=             @������������������������       ��e:59U=              @������������������������       ���
j��<              @                        �=�e?pαe"b[=             @������������������������       �                     �?������������������������       ��"�d�W?=              @                        0]P�?ygvB�=8             L@                         ����?�5�9��=              @������������������������       �                     �?������������������������       �      ��             �?                        ����?�! ��l�=6             K@������������������������       �                     �?        #                 І�s?C�-�S~=5            �J@!       "                 З�Z?�W��]e�=,             F@������������������������       �Ew��E=(             D@������������������������       �`���|Q=             @$       %                 @*��?����[5O=	             "@������������������������       ������J=              @������������������������       ��سݏ�+=             @'       >                 0-3�?ӝ����=)           �r@(       3                 ȃ7z?^y"�[�Q=e            @Y@)       .                  .��?8%-�
O=_            �W@*       -                 ��b�?��;r��'=F            �Q@+       ,                 �=_�?@n/b\u=E            @Q@������������������������       ���Ǌ=D             Q@������������������������       �      @�             �?������������������������       �      0�             �?/       0                 �؉�?��;7�b=             9@������������������������       �                     �?1       2                 0�,�?iڗ���V=             8@������������������������       ��s�a��:=             @������������������������       ��N"��hJ=             5@4       9                 -��?*�[3ǤB=             @5       6                p�s�?l��
5�=             @������������������������       �                     �?7       8                 ��?�/Qf�<              @������������������������       �                     �?������������������������       �      �             �?:       =                  `��? ����%=             @;       <                   ��? mO�J�<              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �??       H                 �\ͥ?TN.v���=�            �h@@       C                 (�e8?�� KǸ�=             @A       B                 ݔ?PX�Z�=              @������������������������       �                     �?������������������������       �                     �?D       G                 �?�V~ju!q=             @E       F                 b?Հ�)�rL=             @������������������������       �                     �?������������������������       ����)��$=              @������������������������       �                     �?I       N                 pN�?���&�%�=�            �g@J       M                 `�ʹ?�Ri�e�=�            `c@K       L                 �X�?#�V���=�            @c@������������������������       �w����|=             3@������������������������       �*�k�<�=�            �`@������������������������       �     ��             �?O       R                 ����?�$�����=#            �A@P       Q                 PUٰ?���פ=             *@������������������������       �����Ij=              @������������������������       ��̑�=             @S       T                 �;X?�\�Fv�@=             6@������������������������       ��'�Q�I=             @������������������������       �2�AK��<             .@�t�b��     h�hhK ��h��R�(KKUKK��h �B�  ׃}�ee>��`��؂��
v dV>ٰ�t�k�߫��r�y�z�	������fY�Կ��TWU������>P���UU忕��HYU�?   iKȲ>�� YU�?  �����>��UU�?%�/|VU�?*A*R�?�>�>��]U�?0�e\�{�>��ݹ���N�JDVU�0�RvUU�UU�&�>0�4XU�?Iܟ�VU�?�fF6��j/��kо����VU�
�E�^U���O�@䗾�:�ZU忥���S����6�V��<��o�ѿe&(CXU�9�>)[{2WU�?~S��UU�?��"?��>��Q4j��Bm�nȋ���m�2�s�����xx��J�UU�|^ZqVU忒���VU�?�(���|��A��TYU�3�&M���0�WU��w��VU�UUMA	ۣ>����1\�>%�1VU�?  ��N{�>lW��UU�?%MӂUU�?UUU����>  芮�>�{VU�?�(YXVU�?�ǰ�VU�?�j#Q_�>ȯ�����>   �*�>lȆpaU�? �V[U�?d=8���>=c��*v�GbHVU忐>%�UU�?�A%XU�?'s6u��>(_��$?�>��+�R��>���s0�ؿ韅���?˩��]U�?<��\��%Zj����l�����?s�5��vSt�9��>`�k
7��?��UU�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K!h�hhK ��h��R�(KK!��h��B8                            @���?;���S$�=�           �}@                        �`>R?`#E5�=�           p}@                        h�[�>���'3��=             7@������������������������       �                     �?                        `�d�?�T� ��=             6@       	                 ��IL?�f�}s�=             4@                         ���?���B�w�=
             $@������������������������       �                     �?������������������������       ���N:��=	             "@
                        �?9?.��_=
             $@������������������������       �T�tV@��=             @������������������������       �l|oW'2J=             @                        ȱ�?�u﨏��=              @������������������������       �                     �?������������������������       �                     �?                        ��U?���XXp�=�            |@                        @Ws�?R"/�.�=             @������������������������       �                     �?                        (d/?Xh֔�;u=             @                        ���m? /�o!=              @������������������������       �                     �?������������������������       �      P:             �?������������������������       �                     �?                        ��LV?��R4n�=�           �{@������������������������       �                     �?                        `("?�X^`_J�=�           �{@                        ��h�>Tr�Ǆ��=%            �B@������������������������       �	��d��=             2@������������������������       ���~�$�=             3@                        `ۭ1?1�?����=�           `y@������������������������       ��h%�{��=             @������������������������       ���c�@�=�           y@������������������������       �     �;             �?�t�bh�hhK ��h��R�(KK!KK��h �B  N���	v�[-g��x��87a��AW|fZU�?W�d��z�� �v��"E&�q>`)CZU��xBK�?���ɏ���'��YU�G���VU�*�*كϾ�uXU�b��\U�mU
_l�����"��>H*�UU�  $��q�>  dH���>R̙�XU�?��YU�?ڧ_\U�?�h����s��.~�]U忥��5p�Ձ)�s	�>���hȿ�O�n��?B��?����I����N��s_�얿@<�
\U�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K-h�hhK ��h��R�(KK-��h��B�	                          �`>R?�ƴ���=�           �}@                        h�[�>N��pI�=             7@������������������������       �                     �?                        `�d�?�T?c͑=             6@       
                 ��IL?Qa,HN�=             4@                         ���?(T�s8�=
             $@������������������������       �                     �?       	                 h��(?h\��Ƅ=	             "@������������������������       �W�Q�<�z=             @������������������������       �[�徒̀=             @                        �?9?`aX=
             $@                        N��S?���RQ{�=             @������������������������       �8p�'�q=             @������������������������       �      p:             �?                        n��W?h�BFkdJ=             @������������������������       � >��=             @������������������������       �                     �?                           �?p�|��~=              @������������������������       �                     �?������������������������       �                     �?                        ��U?��QQ�"�=�           |@                        @Ws�?@�-3퟈=             @������������������������       �                     �?                        (d/?��N`��u=             @                        �j��? �H���<              @������������������������       �                     �?������������������������       �      h:             �?������������������������       �                     �?                        ��LV?���+X'�=�           �{@������������������������       �                     �?       &                 ����?�Mf�=�           �{@        #                 ��{�?����HI�=0            s@!       "                 �U�?Q�;��ȭ=�            @j@������������������������       �0��s��=�             j@������������������������       �     ���             �?$       %                 0*tC?���~���=^            �W@������������������������       ��AI�h!�=)            �D@������������������������       ��7�p�5�=5            �J@'       *                 p祩?Z�EOw�=�            �a@(       )                 �a5�?�BZ��=             (@������������������������       ��2�
�=             @������������������������       ��}�K��{=             @+       ,                  �Q�?����=�             `@������������������������       � 	g��Ĉ=/            �G@������������������������       �Z
�8��=Q            @T@�t�bh�hhK ��h��R�(KK-KK��h �Bh  �(؛QSl>�)��y]�>��WeZU�qn��Q��>*&LT
�>�a��Nl���CZU�?~�l�:��~����J��s�(���?33���>  .�Ě�>"�m�XU�?�%�[U�?  p�T��>�O�0VU�?(ƥsWU�?  ��w1�>L���XU�?�2��\U�?kA�a��C>���u3ľKy�cUU�����ʾA�7ľ�|_�XU���N�XU���U\U忚��h�`>`�(^U�?�M���Q>�=3UӀ�X%���K�>�������?��q�dU�?|�[m,�������ۿJ�a��� �ڼѕ>|ƨ��U�>����n�?c!{��Z���Q�cz�>K��*&¿2��-Y�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K'h�hhK ��h��R�(KK'��h��B�         &                  @���?����v=�           �}@                        ��Q�?�$���v=�           p}@                        0���?q�JA��u=�            z@                        �?g�?�m�j�p=J           �t@                        P!d�?k��B��o=I           �t@                        Ў m?۳�7*l=;           �s@������������������������       �Z
��N�j=           Pq@������������������������       �k\eD�p=&             C@	       
                 ��H�?����N�=             ,@������������������������       �\	O�Jev=             *@������������������������       �      �:             �?������������������������       �      ��             �?                         ���?�@djǂ=X             V@������������������������       �                     �?                        `s5�?c���w=W            �U@                        p팬?�B`��y=#            �A@������������������������       �\KH/M�|=             .@������������������������       ��e17Zhr=             4@                        ��&�?�����s=4             J@������������������������       �$Ӂ!�!c=              @������������������������       ��3~ ��q=2             I@                        ��x�?K %�~=5            �J@                        (��0?����@p=              @������������������������       �                     �?������������������������       �      ��             �?       !                 pg_�?�P"�Ii=3            �I@                        ���?���Zχ=             @                        8��? �d0�=              @������������������������       �                     �?������������������������       �      `:             �?                         8W�?ZL�+[=             @������������������������       ��ܞ><W-=              @������������������������       �)pM�# %=             @"       #                 �Q�?v��lQ�A=,             F@������������������������       �                     �?$       %                 ��ӹ?<�ҭ�5=+            �E@������������������������       ��C��`�)=
             $@������������������������       �����4=!            �@@������������������������       �     ��:             �?�t�bh�hhK ��h��R�(KK'KK��h �B8  �h]�}_>��vpob>U�>8s>����u,X�� �[FF��{-���R>�=��ݲ�ƙ�OC��?&Y�-V��l񆀊ZͿ�$��\U忎
�ZU�/=�S5}�>��+�aU�?��`���>?'�F��>u�����?^�1XU�?�T�e�Zy>F: ]XU�?g�:X�?��a�j��Rq��־~�FW[U���V^U��L���q�Y�|L�����Ȭl;|Ͼ����ZU��ߑhZU忎(Ńx���]p�VU�k�k�UU�?�.|�ѫ�>J*ȉWU�?�0��Qz>�~%�ߖؿd�(�6�?�_h�XU忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KUh�hhK ��h��R�(KKU��h��B�         0                 P�u?�,!'�e�=�           �}@       !                 �C
T?����3��=�             b@                        �U���B���n�=U            @U@                         e	a?�z�a�=#            �A@                        �$?Z?��6w��=             .@                        ���S?�Px�|r=             (@������������������������       �0�O(Se=
             $@������������������������       ���ߗ^�^=              @	       
                 p��3?��b�=             @������������������������       ���f|�k.=              @������������������������       �                     �?                        T�@?�����=             4@                         �Ԧ�?��.qV�=             @������������������������       � �l��_=             @������������������������       � ���<=              @                        �l��?�P}䳛=             .@������������������������       ���!�(��=              @������������������������       �=�	�خ�=             @                        P^N<?妦�xK~=2             I@                        �b'�?u6`T�h=              @@                        �
OW?B7��T=             4@������������������������       �|��"EY=              @������������������������       �Dxg��I=             2@                        ��8?��ح's=             (@������������������������       ����(�"m=
             $@������������������������       �`�<���E=              @                        P^�?�9��M}=             2@                        �5��>Z-vl�=
             $@������������������������       �                     �?������������������������       �jC�*{v=	             "@                          ��~�?�LE��=I=              @������������������������       ��lɶ��5=             @������������������������       ���[OԥD=             @"       /                 �5�t?2�2���=;            �M@#       *                  `���?�}�+.��=:             M@$       '                  �g<�?��9AF��="             A@%       &                  O:�?{���{�=             7@������������������������       ��S)�_�=             3@������������������������       ��#B^}=             @(       )                 ��{�?i&0@��=             &@������������������������       �:g�ͧ0�=              @������������������������       ��e�t=             @+       ,                  ���?Ӈ��v�=             8@������������������������       �                     �?-       .                   ��?c�c��,v=             7@������������������������       �:s�h=             6@������������������������       �      `�             �?������������������������       �      �:             �?1       6                 0Vtv?�3E$��=H           �t@2       3                 H?˵\Q�»=             @������������������������       �                     �?4       5                 p��`? ���{=              @������������������������       �                     �?������������������������       �      @�             �?7       F                 �Z��?꞊�%Y�=E           Pt@8       ?                 �I?��׈d��=,             F@9       <                 @Ws�?j��z��=             7@:       ;                 0a��?R=ˣ �v=             ,@������������������������       ��ɦA;�`=             &@������������������������       �sɛ&��r=             @=       >                 Ш��?|Q�=	             "@������������������������       �l�MV�Ǫ=             @������������������������       �:���}��=              @@       C                 ��>}?��0F�l�=             5@A       B                 ��y?@L_�lS]=             @������������������������       �                     �?������������������������       � xN/�/=              @D       E                 `���?��<�A�=             2@������������������������       �7��θ�=             @������������������������       ����Ly�=             .@G       N                 pG��?�Kp�qA�=           �q@H       K                 ��$�?qv��21�=             .@I       J                 �-�?Bj��J�=             &@������������������������       �                     �?������������������������       �D>F84Y�=
             $@L       M                �J��?e`%���=             @������������������������       �                     �?������������������������       ��_\-�=             @O       R                 0���?�x �%��=
           �p@P       Q                  2V�?��;�
��=             ;@������������������������       �<Yrm9�=             :@������������������������       �                     �?S       T                  �=�?L���+�=�            �m@������������������������       ��k~���=)            �D@������������������������       �z�`n�=�            �h@�t�bh�hhK ��h��R�(KKUKK��h �B�  �n*B�\Z��������>!gǴ�B�����wᬾ�ub�>5�v��k��Ώ��T�ؿ�-$�XU�UU�~̾�>n�XU�?�p��_U�?���f����Ei�y�Ծv�`^U忇�<YU�B���"դ�To*��h�?�� [U忓� �7l�>��2��>�Vq`Ţ>��+�׿����VU�?���:閵>/���WU�?}n�YU�?�E��5���~k����_M��ZU忓�*S`C�V:X�0N��Ţ!VU忰L�[eh�?�b�)�>��b�ˬ>�\$���>�ޕ�W�>1q�w�v�?�o!WU�g	dhϖ�>o�Ej��?ψ$ă�?����K;�><���[U忸Q�S��>��½��?�E�YU忦26_U�?�IW�(���}�%+KѾ}AY�dU�X��]���>�.VU�?[���WU����]y~�IV��C���o�&%CBþ�s�/������PWU�(9)�?����վ���laU�q��k��?׺��N��>��0DK�>��S^U�?���!\U�? �ś��p����῱�����?`k6��0>\��P���>��M��>���\U�T2�Bk��?��ţ���>��d�lU�?�����?U2�?;�9�t�K�����t�ۖѿ��Fi`U忑�u��X�'�<Z��?�ˑ`ǿ�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K]h�hhK ��h��R�(KK]��h��BX         4                 �༡?O���뵟=�           �}@       !                 `���?7��a{�=0            s@                        p�v�?"�S!�n�=�             o@                        �C
T?�������=�            �e@                        �U���*���"P�=H             R@                        ��K�?�t��<Q�=             ?@������������������������       �&�T��ڡ=             <@������������������������       �D�%PtƠ=             @	       
                 �C>?UY�mzv=)            �D@������������������������       �� m�Buc=             <@������������������������       �R�zv|=             *@                        �+?z=x�=e            @Y@                         p��?��1��e�=)            �D@������������������������       �hnaި�=&             C@������������������������       ��'9)��=             @                        @F����E9j�=<             N@������������������������       ��G#���=             :@������������������������       �j<�	���="             A@                        ���s?w�h�=K            �R@                        P���?"�wOD9�=             2@                        �5[h?X&ߴ�=             *@������������������������       ���y8�v=
             $@������������������������       ��LǛ�x=             @                         ��?F��6^��=             @������������������������       �POQ���b=             @������������������������       ��d/��=              @                        �Z��?��XC յ=9            �L@                        @F��h��3�=             4@������������������������       ��:�52�=
             $@������������������������       �SU,L)��=
             $@                         pTF�?
a�M�=%            �B@������������������������       ���o;S��=              @������������������������       ��P֦8h�=             =@"       %                 �-�?<Q
�QA�=8             L@#       $                 ѷz?�k�����=              @������������������������       �                     �?������������������������       �                     �?&       -                  �/�?�$����=6             K@'       *                  z �?�/_uף�=             <@(       )                 ��K?�o9���=             2@������������������������       ���}Y�~=             .@������������������������       ��@ ��j�=             @+       ,                 @�Dv?�U���v=
             $@������������������������       �                     �?������������������������       �n��b^k=	             "@.       1                 P���?�sw��=             :@/       0                    �?����b�=             @������������������������       ��BOjp=             @������������������������       �     �w�             �?2       3                 `���?j�0�'A�=             6@������������������������       �                     �?������������������������       ��	{��!y=             5@5       D                 ���?�o���@�=�             e@6       A                 P%:�?�=k�ݷ�=
             $@7       <                ��X�p?�D�q=              @8       9                  .p�?�c��W\=             @������������������������       �                     �?:       ;                 H!��? �_x7=             @������������������������       � �Mlu}=             @������������������������       �      p:             �?=       >                  �P�? y��gj1=             @������������������������       �                     �??       @                    �?  �N=              @������������������������       �                     �?������������������������       �                     �?B       C                 `��?�7��{A=              @������������������������       �                     �?������������������������       �      0�             �?E       N                  �ŧ?�ӯ76�=�            �c@F       G                 @�?�0�@�"�=             1@������������������������       �                     �?H       K                 �ޥW?#��=             0@I       J                 �?0���=N�=	             "@������������������������       ��P�h�k=             @������������������������       ����,J�`=             @L       M                  ���?�N�E�Jw=             @������������������������       � ��'��=              @������������������������       � 	E�ĕ6=             @O       V                 �/�?�K��=�            �a@P       S                 `Mh�?!�#��K|=!            �@@Q       R                 ����?6��k��q=             *@������������������������       ��P�aEk=             (@������������������������       �      P:             �?T       U                 p�3G?CE<';aw=             4@������������������������       �`�a��wK=              @������������������������       ��8dr=             (@W       Z                    �?!��
�'�=l             [@X       Y                 �S��?�J����=-            �F@������������������������       �7e|XY�=             9@������������������������       ��N��r=             4@[       \                   ��?d�H�W��=?            �O@������������������������       �:�Z&��=#            �A@������������������������       ���8�� u=             <@�t�bh�hhK ��h��R�(KK]KK��h �B�  �)��rH>��ߞ�C~�k�f΋"l>�~k������ 3Ð>k��ȯ>�R���?���]U�?��R3N������1{�x���5�?���d��d�Ӫ�w���q/ooI߿0L L�?��
]R�u>y��5;T�?�0Կ��w��l�>_pf������?��f2j�XU�F���[U�T�D�c~�>���QYU�?����UU��X����>^j����>��	� �?8y�L��?&����x4����H��?3}�ڝǿ}v^�R���[�4�W��3VU�|���lU�z8�����gR������t�����BL���<s�0^U��V��k��Te�	YU�9�?򪰿�V����>t�$։�>�[�[U�?�)"�UU�=�f�����'NZU忞Nq�D)ƿ�ܸF���>���!K�> �����>  ���>?�QJWU�?  ����>�.��YU�?�$(YU�?  ��v|�>o�[U�?  r�0�>Xᰚ[U�?1A;�[U�?lo�!���.P�UU忣b��VU忴��e�;x>�����Ϥ��)\U�?��:6�-��J1ɰ:���'m�YU���v�ҿ]�h�"w�>�7�1XU�?�)6VU��Y)�L��>�+�1_�>ܗ�{�����i*q?r�,XU�PV׼K�>5	&lXU�?SG��,�?�!���b>�iRIQǔ�)@��n⿩p�pV�?Bx���>
�<_���?���p:�ؿ�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K?h�hhK ��h��R�(KK?��h��B�         "                 0�"]?���iZk=�           �}@                        0��?#$@@�n=\           �u@                        �Y&�?nk[�d=           pp@       	                 ��^�?��#�,c=           Pp@                        pִ�?|>:�%k_=�            �n@                        p ��?��F���\=�            `n@������������������������       �IF��3�Y=�            @k@������������������������       �����`=             9@������������������������       �     ���             �?
                        |�L?i\�:+�|=             1@                        P���?
�3��=              @������������������������       ��|�V�~:=             @������������������������       �      p�             �?                         �{��?P~�D�7L=	             "@������������������������       �DuXjܼ;=              @������������������������       �       �             �?                       �o|?�x3�\F=              @������������������������       �                     �?������������������������       �      `:             �?                        �ˤ?pol{n�}=U            @U@������������������������       �                     �?                        PeT�?=vlp��x=T             U@                        @?,�?��I�T�}=             6@������������������������       �                     �?                        0kz�?{�H-�r=             5@������������������������       ��ĥ��Mu=             @������������������������       ���J��g=             1@                        @��8?���|�t=>             O@                        @*t3?�@�F�t=,             F@������������������������       ���f=+            �E@������������������������       �      ��             �?        !                  u�?gG� �j=             2@������������������������       �(F�lY=             1@������������������������       �      p�             �?#       &                 p�]?�Y�yaa=|             _@$       %                  p��?U��E0^�=              @������������������������       �                     �?������������������������       �     XH:             �?'       6                 �#=�?!�֢Z=z            �^@(       /                  ����?՞���X=5            �J@)       ,                  ~?��ۻh�C=             3@*       +                 Pl?ֳ��)==             &@������������������������       ����⋛+=              @������������������������       ��O��"'=             @-       .                 ����?��/aS�0=              @������������������������       �,� e���<             @������������������������       �                     �?0       3                   ��?P���\="             A@1       2                 ���?h�Yx�He=              @������������������������       �                     �?������������������������       �                     �?4       5                 �uU�?޵E���G=              @@������������������������       �E��/X8=             <@������������������������       ��3"c=             @7       8                 @sߦ?C��5,Z=E            @Q@������������������������       �                     �?9       <                    �?��1REV=D             Q@:       ;                 ���?�i�%=             >@������������������������       ��f��5=             @������������������������       �N��x=             8@=       >                 �N��?B�f�N�a=&             C@������������������������       �.J5!m=
             $@������������������������       �t���:!W=             <@�t�bh�hhK ��h��R�(KK?KK��h �B�  ��]��GL><��`��\���yIEv��;�|q��U�Y{�j]�t��~�j=f5ſ�e@WU�����YU�?^�~CVK�>  ��9�>�ֈ�VU�?6P_3\U�?�O��rw���d:VU快�TLVU�?���4B�ž��5lXU����YU�P��)��>����\U�?#�V��v>�� g���>3��[U�?�q���>i�80��?ke΍���?�s�2AA~��Az�t>�p�Ԓ���cA1\U�?�	�~J��� ��J!���YU�Dd�гԀ>  �Cy��>y �ZU�?��~[UU�?-�0Ԗdy>V��z6�>M��S�c��-�
����[bD��տ���KVU�  8,��>��.�UU�?�ٲ�VU�?����ɩ�>   "�>�&TWU�?SG�YU�?�T?��>He����?��@%�-�?�ѐ:��S���/XU忲���{H>��Φ���>�� VU�?��f�UU�?=�5�z���d�vO�<���?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KGh�hhK ��h��R�(KKG��h��B�                             ҏ�?+���r��=�           �}@                        �7~�?C��E-�==            �N@                        �w4�?���Ԁ=<             N@                        ���?��O|���=)            �D@                          ���?s˽E�{{=#            �A@                        PeT�?*z��x=              @@������������������������       ���1��n=             8@������������������������       ��"9s��=              @	       
                 p��?����w=             @������������������������       �d�.D!�B=              @������������������������       �                     �?                        �;�j?�/Q���~=             @                         `���?Xm�@�s\=              @������������������������       �                     �?������������������������       �      �             �?                        p8��?����D=             @������������������������       �  &Z��<             @������������������������       �      |�             �?                        0o=�?/�gI�w=             3@                        ��O�?�F�UM�=             @������������������������       �                     �?                        `E��? �!�W�<              @������������������������       �                     �?������������������������       �      �             �?                        (�3?��6
[U=             0@                        �9.�?g8GkDXe=             @������������������������       �                     �?������������������������       �rr/�A3=              @                        P7&E?N��bV@=             *@������������������������       �                     �?������������������������       ��2U�:�&=             (@������������������������       �      ��             �?!       <                  ����?٧�M�ށ=�           �y@"       1                 ����?r�T�-%�=�            @l@#       *                  v_�?���>��=�            `h@$       '                 ���?���=�            �e@%       &                 ��h�?����߈�=�            �c@������������������������       ��Ir5ǃ=�            �a@������������������������       ��
ԯ �=             1@(       )                 `7h�?��t�%�r=             .@������������������������       ���0�aq=              @������������������������       �}��P-gW=             @+       .                  t0�?M�[���=             6@,       -                 ��?J��ǅ�=              @������������������������       �                     �?������������������������       �                     �?/       0                ���K�?pb��O>�=             4@������������������������       ��i	��4�=             @������������������������       ���v�^T=             ,@2       7                  ���?4���/�=             ?@3       4                 `��?�M�S�o=             :@������������������������       �                     �?5       6                 �P�?B͜�Vxg=             9@������������������������       �V�Cq�(r=
             $@������������������������       �5_���iQ=             .@8       ;                 ���?�˘�≚=             @9       :                 ��o?r*P��<             @������������������������       �                     �?������������������������       �SG�k:<             @������������������������       �                     �?=       >                 ��1?�<�B��g=�             g@������������������������       �                     �??       F                  @���?J��F��f=�             g@@       C                 ��'�?wʬ�Vf=�            �f@A       B                 ��{�?r����d='            �C@������������������������       �1y�5�^="             A@������������������������       �NVdX?p=             @D       E                  �6�?�r���e=�             b@������������������������       �������y=              @������������������������       �:q反b=�            �a@������������������������       �      �:             �?�t�bh�hhK ��h��R�(KKGKK��h �B8  E4
��$e�x�*:s��Ft�f����)=�ʍ���O�u��h W��ؐ�&�cԍ�[?�Yȹ�޿]M>ΚE����VU���9�YU��t>ๅ¾� ������%�VU��`��UU�?F��P��ɾt���YU��缲XU忾:����r>����3�>~��[U�?  [�^�>-��UU�?F�VU�?��������!�tE���ºXU忡#�VU�D�!��|�Sx$�VU�?����UU��l�^U忛���v(a>�mA�S��>�&�r���>F|��2ʅ>� `�h�>��%峛�?GK�2�?B˯䝘��5}[5XU���9�iլ��Q�w�>  ��B�>��XU�?�P�dU�?%�TP��>��n��5�?�Y�/���*�Z�c���`1;����<
ܽYU���FnH�����0XU��NV ú�ڷ�:f�>'�j�nJ�1b�dUU忧�SVUU忮u��]U�?�CVV������YU�*�L̂��3�v���sj�vDJ|>O�e.�������E��?�vqBe��Q�ZU�"C��s-ֿ|��WU�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KAh�hhK ��h��R�(KKA��h��B8                            ҏ�?�K����=�           �}@                        �7~�?O�q���==            �N@       
                 ��k�?| _�B�=<             N@       	                 ����?��7���~=!            �@@                        ���?�~~>@pt=              @@                        0B��?�N��.�o=             ?@������������������������       �������o=             7@������������������������       ���M��X=              @������������������������       �      ��             �?������������������������       �      �:             �?                        X��?�wx��z�=             ;@������������������������       �                     �?                        �Z�?�z�y|�{=             :@                        Pi��?���x�=             ,@������������������������       �ѝ-�fJl=             @������������������������       �輒��w{=             @                        0.��?N*�vV=             (@������������������������       ��I�T�K=             @������������������������       ���=>�<=             @������������������������       �      ��             �?       0                  ����?��o�k��=�           �y@       #                   ���?~
G���=�            @l@                        `@��?�M��ֆ=�            @g@                        �j[?����Ry�=�             d@                        `}��?��M�e�=M            @S@������������������������       �X���Z�=K            �R@������������������������       ����g�x=              @                        @l�?T�%��8}=T             U@������������������������       �W�AX�|=B            �P@������������������������       �xt�2v=             2@                         `��?����A�}=             9@������������������������       �                     �?!       "                 0�2�?�@o�t=             8@������������������������       �*�w��;=	             "@������������������������       �3��)\zz=             .@$       +                 �؉�?+���_��=(             D@%       (                 @Ws�?��]�N�=$             B@&       '                  L��?�x:�=             &@������������������������       ����#�t=
             $@������������������������       �      p�             �?)       *                 P�p�?�'y�y=             9@������������������������       ��o�-�<�=              @������������������������       �~�ӛ�Uj=             1@,       -                 �v��?�q�����=             @������������������������       �                     �?.       /                  ���?T�

�g�=             @������������������������       ��P7ylU=              @������������������������       �      p�             �?1       2                 ��1?�F���Mr=�             g@������������������������       �                     �?3       :                  ��?�!3�R�q=�             g@4       7                 Ш��?���i�k=}            @_@5       6                 0�2�?#��[Yj=V            �U@������������������������       ���&,��g=U            @U@������������������������       �      �:             �?8       9                  �!�?����)m='            �C@������������������������       ��d�	��k=             :@������������������������       �}�}o�0e=             *@;       >                 p�,p?q�yx=;            �M@<       =                  $��?��Rq�=             5@������������������������       �b�LQ~��=	             "@������������������������       ��6�uit=             (@?       @                   �0�?~_tR�gM=&             C@������������������������       �hC�y��h=              @������������������������       �>ń�D=$             B@�t�bh�hhK ��h��R�(KKAKK��h �B  X�I]tW>.	\r�>̧�y�A�>��Hه>̻��X�>@B��:��>�2+����?"�8�y3߿t���YU�?6��][U忩D�<q�>~��W[U�?;�>�
���ܴ>e���ީ�?C�\XYU�?�o���`>
�pk}�?7f�CVU�iי�^U�?�5p�o�H���Q��r��W�_����+Z�a����&����X�+�dʿ��I�YU��U�E��V>����?�?B3%��ڿF�(Ǚ�>Ag�
[U�?���)�*�>�:$���࿙o��s��?�X�d�K(H�|����;�$�>�س���?��ZU�?c��HK��R����<���Ͽ��X̂�о=,�pcU�Y*\�����ΚWU忚��[U忼�_k�݁>V�YU�?�5[���>׭��7���n|w>�R��5�?���=YU�?�S��8F����{�x�ٿJW��*��?�����>��JA��>R�'��'�?<��Aΐ�?�`do��c>������?Wj묛���t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KEh�hhK ��h��R�(KKE��h��B         0                 �)�?���ȠbR=�           �}@                        @�_�?b��lnoR=�           �|@                        ��ð?!0��)�R=�           �y@                        ��\�?g���kQ=�           `y@                        ���?��'&=�C=�            `o@                        �6J�?�E�*-B=�             n@������������������������       �}`(%ܳA=�            �m@������������������������       ���@�<0=              @	       
                 ��d?L��wL�P=             &@������������������������       � ����P=             @������������������������       ���8��=             @                        zL&?�$�}�\=�            `c@������������������������       �                     �?                        ��ؿ?��PVw�[=�            @c@������������������������       ��yM��?s=             *@������������������������       ���~r�U=�            �a@                       ��&��?�/�5��=              @������������������������       �                     �?������������������������       �                     �?       #                 �.KR?�e7���N=3            �I@                         c
8?2��݀�]=             *@                           �?�4l�?=             @                        @��?K� ���J=              @������������������������       �                     �?������������������������       �     ��9             �?                        `�@�?@���s� =             @������������������������       ��e��Ī�<             @������������������������       �                     �?                         PUٰ?H���_=             @                        `��?D��ml�!=             @������������������������       � ȟ���<              @������������������������       � �j��0�<              @!       "                 T��?�7�i.=              @������������������������       �                     �?������������������������       �                     �?$       )                    �?�f-�-@>=&             C@%       &                 ��Oa?�ǒ;��=             *@������������������������       �                     �?'       (                 p��?t�� ��=             (@������������������������       ����+"�=             @������������������������       ���_k���<             @*       -                  �j�?��&e�B=             9@+       ,                 `���?9L���G=             (@������������������������       �u�\)4�2=              @������������������������       �8� o�;=             @.       /                 �;X?�8h�O==             *@������������������������       ��xܸ�i=             @������������������������       �����s�<
             $@1       6                 p�ռ?�VEk��E=             *@2       5                  ���?`�=�^1=             @3       4                 ؾ��? :2!5��<              @������������������������       �                     �?������������������������       �       �             �?������������������������       �      0�             �?7       >                 ��?�	<-=
             $@8       =                ��}r�?���%=             @9       <                 �D�澠5,:��<             @:       ;                  �9��? �d��#�<              @������������������������       �                     �?������������������������       �      :             �?������������������������       �       �             �?������������������������       �     �:             �??       D                 �/��?�wcс��<             @@       C                �qd�?�{��i�<             @A       B                 �)�(?���n�.�<              @������������������������       �                     �?������������������������       �      ��             �?������������������������       ��T��O5�<             @������������������������       �                     �?�t�bh�hhK ��h��R�(KKEKK��h �B(  ��8���R>��0�	�D>�-a���_>��Rp��X>l�)}[�bEB32:���[L�]���RjVU忰Y�������V�VU�VV�UU忤
�8�9{>�~�WU�?T�gG�2x>�89
�)�?Pz5����?�
OyL��>�i�VUU�E}YYU�?��5E�:��`M��r���Y�z�x��9�]���Q�~VU�烙cUU�?��:F�^>��uUU�*��UU�?[Pp�]���6W8�S��w�,VU忣�%�UU�.���㽾�Y9�WU�˻�%XU�4	LEi��N�6�y~>��VU�?��J�NMu>��UU�?���[UU�?���	؆�����ڟ�����Jڿ�̙VU忞؉�r�s>�4�UU�?^��qUU�?[;���>  ���{�>  �s��>��tEVU�?�j?^VU�?D-�WU�?��v>>��>  �Af��>  ��͞>  �AX�>�.��UU�?���VU�?\l_�UU�?c��_UU�?D����\��4���/�F����a����[UU忤�fUU��b�_UU�?���UU忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K_h�hhK ��h��R�(KK_��h��B�         *                 )DW?;o�#ݨp=�           �}@                        ���p?:�ͱ�:t=b            �X@                        @�p?�f+�?~=-            �F@                        0�G?���	}�{=,             F@                        �j�a?tҙ0ր=             >@                        ���U?�����hq=             6@������������������������       �5�E�sz\=             *@������������������������       ����B�z=	             "@	       
                  �G�>��u���=              @������������������������       ����{�x=             @������������������������       ���`A�WU=             @                        0��o?Tu%�\]=             ,@                        ��?>�B�%U=             *@������������������������       ��Mq�W�M=             &@������������������������       ���H [�;=              @������������������������       �      P:             �?������������������������       �      �:             �?                        PeT�?jx޹ѵd=5            �J@                        ��?���d=*             E@                        @F�����7La=%            �B@                         `�J�?�zԶ:�[=!            �@@������������������������       �
̹�;9t=              @������������������������       �LXf��S=             ?@                        p��N?z&����i=             @������������������������       � @P��J<              @������������������������       � �w1Ȓ3=              @                        �t�E?�F\��Y=             @                        �l��?���8�L%=             @������������������������       �      @:             �?������������������������       � ��
=             @������������������������       �     �V:             �?        %                 �vs?l����|\=             &@!       $                 ��1i?���ZR=             @"       #                 �;A?ֳ�%�;=             @������������������������       ���� �3=             @������������������������       �      �             �?������������������������       �      0�             �?&       '                 ��? xj\��%=             @������������������������       �                     �?(       )                    �? �e��<             @������������������������       �                     �?������������������������       � PJ��<              @+       J                 вeh?l	1j�>o=v           `w@,       ;                 �?o�?0��ԚZq=�            �b@-       4                 �N��?�.6��z=@             P@.       1                  T?�X4��j=0             H@/       0                  �\�?�66�zf=+            �E@������������������������       ����,ke=	             "@������������������������       ��()��c="             A@2       3                 P��n?~�B8.�r=             @������������������������       ���<��BR=             @������������������������       �                     �?5       8                 P���?�����=             0@6       7                  @?��?�)XΈ|�=              @������������������������       ���ҚV�!=              @������������������������       ���C�>�u=             @9       :                 p��A?����zt=              @������������������������       ����Ә[f=             @������������������������       �      P�             �?<       C                  �P��?:.3N>fb=U            @U@=       @                  �7�?*�Hb�k=             :@>       ?                 �༡?-�>$Uf=             7@������������������������       �P�[o=             &@������������������������       ��#&!|E=             (@A       B                 08��?c���u=             @������������������������       �                     �?������������������������       �J�$u�6=              @D       G                 �2z�?�Фu�JY=;            �M@E       F                 ��r�?O�q�K�W=             &@������������������������       ����T��,=              @������������������������       �����x8=             @H       I                  �p�?=��J�EW=0             H@������������������������       ��z>R�Ec=
             $@������������������������       ���[O�E=&             C@K       T                 pc\�?��,�l=�             l@L       M                 Pa�l?��B׷p=:             M@������������������������       �                     �?N       Q                 �7\?�4I��ql=9            �L@O       P                 �FX?���Kq=)            �D@������������������������       ���䄿n=(             D@������������������������       �      �:             �?R       S                 ��c?JU[c�;=             0@������������������������       �                     �?������������������������       ���JM2=             .@U       X                 Pf�b?�o�v��h=�            �d@V       W                 �m��?�����G�=              @������������������������       �                     �?������������������������       �                     �?Y       \                  �~��?iW����d=�            �d@Z       [                 Ć?n��b(3f=3            �I@������������������������       �B$�E�t=	             "@������������������������       �atY�SW=*             E@]       ^                 �Ò=?�8W��<c=r            �\@������������������������       �Q��V".v=             ;@������������������������       ���i��	S=W            �U@�t�bh�hhK ��h��R�(KK_KK��h �B�  ��o3�\��"��*N|>6�
}�j� �� �k���r˩Γ��רX�f�>��R�=�����e|��?�}5�T������YU��;�ɥ�Y�yG1��>9f�Ѫ�>H��VU�?j��<VU忽7��WU�?��YU�H@����>^�cɕ��>z��8�"�>Ҕd��،>��H��޿u��v^�?  �.~а>����UU�?���WU�?��\$�Ҵ>  (W��>�]�WU�?6΅YWU�?���pUU�?_M>aԄ��2��I�>��T��`>w��UU�?ß�4VU��[FWU�?i��=B��3�q�UU�|�2��k�1�VU�;��VU�s�{>߃p��
����_�z�Pu���[����pC����
�na,k�?�)�ۿ2y`��>���
9��?o���XU�?��5
J��ԯ7��þ��>VU��^�ZU忰�>�%Rs>�G�{v?ʿ[�QXU�?92��b���Z�M�>�<�p���>����;��?��ߍj��A�)Xs�>{h`�XU�?��5��4�?!4��s���,��`��>^zVU�0��VU�?�����؏���akWU�	,a�RpϿ�O��5c>#1�̗>k���YU�?LYz΂J�>$?^��G�>tFA��?��YU�?�J?�L��zF�VU�ߖDEVU�!t�3�k�1�Ǿ�+�CWU心��K[U��i҇�[f�-�h�����:�]XU忞,�u:G����[�r7h>��8f�e�?]�+};"п�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KKh�hhK ��h��R�(KKK��h��Bh                          ���p?Fht!�sr=�           �}@                        @�p?�83o���=M            @S@                        0��?�S���~=K            �R@                         !��?; ��Y�{=F            �Q@                        ���r?���&�Cy=E            @Q@                        �"b?$FH{�y=>             O@������������������������       ��NT
�Qz=3            �I@������������������������       ��g잩h=             &@	       
                  �Z�?ĵ�K�X=             @������������������������       � 'ΰdI;=             @������������������������       �7�b�2=             @������������������������       �      ��             �?                             ��`���=             @������������������������       �                     �?                        p�q?�y���`=             @                           �?�RD=             @������������������������       � ^��q�<              @������������������������       �      :             �?������������������������       �                     �?                           �?`3�V`D_=              @������������������������       �                     �?������������������������       �                     �?       ,                 �?�7���m=�           �x@       %                 x��?�޳=�f=#            �A@                         @F����7�b=             ?@                         `���?�2�� ]=             <@                        `7p.?yøB�t=              @������������������������       �                     �?������������������������       �                     �?                        @*tC?�\�zT=             :@������������������������       ���q���O=             4@������������������������       �L�����N=             @!       $                 ���?�U$���f=             @"       #                  pS��? P{��>=              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �9             �?&       '                 �4k?����<$=             @������������������������       �                     �?(       +                   ��? �ݲ��=             @)       *                 Њ�(? xJլ��<              @������������������������       �                     �?������������������������       �                     �?������������������������       �      T�             �?-       <                  �~��?��Sv(�m=h           �v@.       5                  �P��?)9��t=            �_@/       2                   �G�?�JmXh5b=Z            �V@0       1                 �7~�?�D����Y=(             D@������������������������       ��Xی>�U='            �C@������������������������       �      @�             �?3       4                 �J�?%wF��d=2             I@������������������������       ��tsFڂf=             9@������������������������       �-GҌ�[=             9@6       9                 �Y�b?]����Ѕ=%            �B@7       8                 @�C�?��푗�=             0@������������������������       ����B;�=             @������������������������       �<g��~=             &@:       ;                 �ҍw?z%��=             5@������������������������       �                     �?������������������������       ��Q�B�y=             4@=       D                   �P�?&L��dh=�             m@>       A                 ��ܳ?~޸��v=             (@?       @                 ����?9C��w=              @������������������������       �|��K�h=             @������������������������       ��1v��Si=             @B       C                 Ш��?���BQ=             @������������������������       ��sw�|�=             @������������������������       �                     �?E       H                 ��I�?0؜~uXf=�            �k@F       G                 �(+�?�ɑ��n=.             G@������������������������       ����o�k=             :@������������������������       �TW��|*g=             4@I       J                 Pֵ?��C$s�c=�            �e@������������������������       �s�1MI�p=             :@������������������������       ���t%3`=�            �b@�t�bh�hhK ��h��R�(KKKKK��h �BX  B�kdS>L���	�>�S
���x>�H�Q�O>��t u�p>�]�`Qt�><ZS�p�?�S���?Ye�ZԬ�FxtWU忆Oi#VU��S��YU忾��
�>zըP[U�?��HS�4�>�'�0=d>.�[�UU�?��VU忔+�[WU�?  D̥k�>���[U�?ƒ]�YU�?��^	�O�MH2O�:��t@e�s���gT�ʤ��bT�^�H�>�|'�UU��}��WU�?!;��A*���"����߿\d(���?o�.�����z�G?й��mK~ZWU�gWzDXU�fV�UU�fI����n@��WU���׷���+�Ӹ���jyWU�$��TWU�e��'WU志�u��aW>o�G�%�>f��kϽ�=@#�d���>=q�����?�M�WU�?��p�����e�mڿ3�����?�[���m�>uQ�Аy�>�E�nZU�?�� 7���?��8�܃>���YU忑��wXG�?4v�g�wό��6���|�#>���J���ӿ��Y�XU�hp&��O�>U���UU�����VU�?d/'��M�SioAq�>�R��8D�?O�g�Ͽmݳ�r����pvڿ�<=y?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KIh�hhK ��h��R�(KKI��h��B�         0                   p��?��X6E=�           �}@                        �6Sz?����C=�           �z@                        @8��?k���ZSF=[           �u@       	                 ��K�?�s�gE=Y           �u@                        �3��?#�E���O=�            �`@                         �/�?tå���M=�            ``@������������������������       ��@?�w�H=|             _@������������������������       ���0g�e=             @������������������������       �      P:             �?
                        @�P�?��6"==�            �j@                        ��?�z�3�D<=�             i@������������������������       �pvǳQ4=�            �c@������������������������       �ϣ�v��H=,             F@                        ��X�?�|w�(M-=             *@������������������������       �P�]me�'=             @������������������������       ���D� @=             @                        @���?>,�c��j=              @������������������������       �                     �?������������������������       �      /�             �?       #                 @EE�?��g�z0=Q            @T@                        P���?n���W(=<             N@                        ����?ě�FwE(=,             F@                         ��d�?>�O�82=             ?@������������������������       ��(V8&�!=             &@������������������������       ���Z��<             4@                           �?ӟ�С23=             *@������������������������       �|p���E�<             @������������������������       ��B�-=             @                         @L��?Fx9�	=             0@                           �?d��v=             @������������������������       � B0���n<              @������������������������       �������<              @!       "                 ���?p��z�<             (@������������������������       �  �/�w
<              @������������������������       �:�`U�إ<
             $@$       )                 Pα�?7��i7=             5@%       (                 ����?&�z�S�P=             @&       '                 ����?�@0���5=             @������������������������       �                     �?������������������������       �@�d����<             @������������������������       �                     �?*       -                  ��?�^`��<             0@+       ,                 ��?�#.����<             @������������������������       �n����f�<             @������������������������       �      �9             �?.       /                 @;;�?�Y�Ļ�<             &@������������������������       �                     �?������������������������       ��ȕ��<
             $@1       H                 �2*�?֔����M=,             F@2       ?                 ��=?¦����A=+            �E@3       8                 0�H�?!�2�2=             6@4       7                  �2�?��kw��0=             (@5       6                 �c��?�ŕrH]'=
             $@������������������������       ��jW�)�=	             "@������������������������       �      :             �?������������������������       �  ���8<              @9       <                 `5�?� � �=
             $@:       ;                 X��?@��w�F=              @������������������������       �                     �?������������������������       �                     �?=       >                 �GD�?5?Z��<              @������������������������       ��z�B�<             @������������������������       ����O�<             @@       A                 9�H!?�J���F=             5@������������������������       �                     �?B       E                 p�;_?���*�==             4@C       D                  �{��?�1E
�P=             @������������������������       �0��ɏ.V=              @������������������������       �51z�&�=             @F       G                 �m�?L���)=             ,@������������������������       �                     �?������������������������       �>�ĭ%�<             *@������������������������       �      t�             �?�t�bh�hhK ��h��R�(KKIKK��h �BH  �T�Ӑ�B>�׫���1��|XZ��"���^��  ��~[>��w�B�c>;N��Ǣ?�2���?�<MWU�lB D��p������u�����y'̿F�/�߿��pi��>��8VU�?Tx�W��?��?V_�>g�1�WU�?Oޔ�UU����sGv>5FGm�>����zl�>t�y��$�>�P��UU�?����UU�?;�Y�>gV��UU�?�x0VU�?�Ņ1I�X���B�\\��&!�XUU�?"YF�UU�   t@�R>�0)jUU�?t�z^UU�?�� �
rg�P������f�]{���%VU忠� nUU�?��m�VU�  @~�e>�� ��x>�h�sUU�?�$\�UU�?   R>�04kUU�?�:�]UU�?	;@�� �>����8x>��C�"b��ft�=煾�����x���E�UU���k�UU�?�7VU�fff(�O�>  �����>3���UU�?&K�VU�?   g?*j>b�]UU�?��~UU�?I0ϕ}��>m�H*WU�?N��4�:�>�	�X���>��WU�?x
�P3=�?���Aq>yD;�UU�?;��6���?���7XU�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KYh�hhK ��h��R�(KKY��h��Bx         2                  (w�?�(P}wW=�           �}@                        �/��?�L�GJ�Z=T           @u@                        ��P�?0/Vt�Z=A           t@                        _��>Ha9M�\=           �p@                        �0?#?�2��yg=             3@                        P���>��j���5=             @������������������������       �!�Jr��=             @������������������������       �                     �?	       
                 ��_0?b�NP�m=             (@������������������������       �                     �?������������������������       ��Y�h�Z=             &@                        ���>�y�[=�            �o@������������������������       �                     �?                        P���?�{&v\�Z=�            `o@������������������������       ��BGkCZ=�            �n@������������������������       ��t����X=             @                        p��?��pC�mM=2             I@                        ��Z�?u��"�XS=              @                        �@�w?@���Aw=             @������������������������       ��g�L�<             @������������������������       �      0�             �?                           �?��ّ��K=             @������������������������       �3Нp�+=              @������������������������       ��Y8h=�"=              @                        H~��?x���E=*             E@                        ��{�?�}��HhI=             4@������������������������       �Hn���1=             .@������������������������       ��{����N=             @                         ���?D�m9�9=             6@������������������������       � �J��<              @������������������������       �J��ʑ�5=             4@        +                 �I��?�"fwU=             3@!       $                 \��X?j�	CE=             .@"       #                  ��n?��zC�X=             @������������������������       �   ����;              @������������������������       �     `�9             �?%       (                 ���~?g���'dB=             (@&       '                  �JV�?�:q��&=              @������������������������       �                     �?������������������������       �                     �?)       *                 Dm�p?DH�5��9=
             $@������������������������       ��ŎFߌ<=             @������������������������       ��֝��<             @,       /                  ���?m50�"d=             @-       .                    �?`��t(=              @������������������������       �                     �?������������������������       �      �             �?0       1                 �K��?`�<(��;=              @������������������������       �                     �?������������������������       �      0:             �?3       H                 �H�9?W�΅�QK=�            �`@4       ;                 �I�?x����IV=4             J@5       :                 ���?ɷ�N��Y=             >@6       7                 ��=�?��5v#ZP=             =@������������������������       �                     �?8       9                  �Q�?�����H=             <@������������������������       �S���>=              @������������������������       ��O�?=             4@������������������������       �      p:             �?<       C                  0�?rXF-5=             6@=       @                 @��?6���8uA=             @>       ?                  �_�? �����<              @������������������������       �                     �?������������������������       �                     �?A       B                 ��N�?Z`�9�{)=              @������������������������       �                     �?������������������������       �    8��9             �?D       G                  �6�?V9�&=�<             2@E       F                 �*8�?X�q����<              @������������������������       ���k6��<             @������������������������       �-d�n�O�<             @������������������������       �yk���n<
             $@I       L                 `�C?:�``9=P             T@J       K                 �8��?�O����$=              @������������������������       �                     �?������������������������       �                     �?M       R                 `�4x?���=N            �S@N       Q                 w?μ_�?�+=             :@O       P                 �1�?3n�)��$=             9@������������������������       �"��c��<             .@������������������������       �	o5IW5=
             $@������������������������       �                     �?S       V                 �p�?�w�JQm�<4             J@T       U                 �,U�?��ܫ��<,             F@������������������������       ��q� 2��<             ,@������������������������       ��T��sLZ<             >@W       X                 @���?���Ծ=              @������������������������       �                     �?������������������������       �͙e��;             @�t�bh�hhK ��h��R�(KKYKK��h �B�  �)��R������Q>Jc����=Bv�HS$`>a_���R����~�n��>4��J�?ĝ�vVU�?C�MC���/qEYU�X|��~�ֿ�F_C4k>�b<mWU�?�* �$h>�:
z�p�?�Fc%R�?����х�&�_�����U���������VU�IuKWU忊�<g��u�_���?�)�BVU�-1�:�st��(e��xfJ�ϿG!^�VU�l��;,�g>�/��UU��>�ԪL�?�������>��⾅>	���'y���&Y�UU�;9�\UU��uɗ��>  Xw+H�>�C%VU�?�wުVU�?����F�>���9VU�?QQ��UU忬��Kx�>�:��u>#Y>�UU�?�f�UU�  �(9�>MO��WU�?�Oz�VU�?L�bƂ{��n�����!<�Dt5�� ���Q���TF�WU�`5�|o|��R�+�zQ�?�WK����j��XU�t��/D[p>��n6͡>  h��z�>��,�VU�?�:VU�?�$Ԋ�~�>�lx�UU�?b�UUU忺����Og�[{ru"*y�����UU��N�jUU�R��WUU���)n;4�  8�a�>EsoXWU�?�9��WU�?c�ǝi�$�C�~�o�ž��w����oUU��
",VU��|�NVU���U���M�f��L��>�����UU�z1�WUU�ߍ@�G�k� %I�UU忝�oUUU忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K9h�hhK ��h��R�(KK9��h��Bx                          _��>�J?���[=�           �}@                        �0?#?���<h=             3@                        P���>�5㎱&6=             @       	                 �>W�>g�Ow3=             @                        ��ڢ>0�6���=             @������������������������       �                     �?                        �]/%?0sr��<             @������������������������       ���6a�^�<              @������������������������       �                     �?
                        0�!�?/2�v5��<              @������������������������       �                     �?������������������������       �      �9             �?������������������������       �                     �?                        ��_0?��ǋ�yn=             (@������������������������       �                     �?                        ��E?�5���[=             &@                         �vg?(8yNH"U=             @                        ����>�ޫ �@=              @������������������������       �                     �?������������������������       �       :             �?������������������������       �                     �?                        xQ�X?��ftN=              @                        X[cp?#��3�>=             @������������������������       ��v�YE�<             @������������������������       �n�rW�!=             @������������������������       �                     �?                        ���>bG��(�Z=�           P|@������������������������       �                     �?       ,                 ����?l��m|VZ=�           @|@       %                 p�!�?�	��]=8           �s@       "                  ��?0m�8�\=�            �`@        !                 �C[?ip�T.a=             .@������������������������       �                     �?������������������������       �_����]=             ,@#       $                 `[�?���A�Y=w            �]@������������������������       �ƛq8��W=o            �[@������������������������       �\���W=              @&       )                 _5?��O�]=�            @f@'       (                 ���?:p �@KY=W            �U@������������������������       �62�,W=V            �U@������������������������       �      `:             �?*       +                 �<�?�2Z�`=[            �V@������������������������       �xv��/a=              @@������������������������       ���.���[=;            �M@-       2                 �D���o��vR=�            �a@.       /                 ����?nZ�-�`=1            �H@������������������������       �                     �?0       1                 �I�?�|��q[=0             H@������������������������       �݅j�fc=             :@������������������������       ���>���/=             6@3       6                 `�C?Uzv�աA=[            �V@4       5                 �H�9?�X���X=             @������������������������       �aο�c0@=             @������������������������       � ���<              @7       8                 `�4x?,��P2_7=T             U@������������������������       �.����E=             >@������������������������       �5��P�#=6             K@�t�bh�hhK ��h��R�(KK9KK��h �B�  �=X�18B>������>�,�]��1�q���s���5���	ܿ�UU��}l;$z�w�kUU忝!L�UU�_��>-n>�/�UU�?�:�YUU���uVU��z!}6`�>�p�XYU�?b:�e�>��:C-�>  p�2�>a�VVU�?� ��UU�?,��WU�?�a�e�p>+ڴ8d�r��e��UU�?�s��UU�_O��VU�?I)E5"�A/bWU�8�MF>4Ѵ�)Cd��j�l|f>5S��-���@!SVU�?��7Yj�促a)rV_{>g����Ķ?���Gˋ�?BX���8z�O\QR�����Ku(��ӿ�'�nWU�?��۸<;>�z�B9�?�����ſ�G��w>ex��(�>gB�XU�?lY�}<t�>�h���'�?@-C���ҿ8��]p3'�V��#����3e�Lֿ�Cw3WU忟|���4e>ƞ9 ��?��]?���t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K1h�hhK ��h��R�(KK1��h��B�
                          �\�?'��R6=�           �}@                        �$��?��k�e=�            @j@                        0��?��3o3=�            @i@                         U�?���m;O=�             i@                        ��?vK恘�=�            �h@                        �e�?�	Pt�<�             g@������������������������       ���EsO�<�            @d@������������������������       �e7t$"=             7@	       
                 �J�?1����z4=             ,@������������������������       �                     �?������������������������       �禥w_#=             *@                        ����?��kVC=              @������������������������       �                     �?������������������������       �                     �?������������������������       �      l:             �?                        `|)�?�Xf��)=              @                        �N��?�zW�U�'=             @                        C�? �,,���<              @������������������������       �                     �?������������������������       �      �             �?������������������������       �      �9             �?                        �rn?�X�s��<             @������������������������       �                     �?                        �&+�?n���<             @������������������������       ��i��z<             @������������������������       �      p�             �?                         �D��?���}~A=           `p@                        ��)�?�E��f=             @                        ��j?֘0Vb�5=              @������������������������       �                     �?������������������������       �                     �?������������������������       �      @�             �?!       "                 �aH�>Vw��-N?=           0p@������������������������       �                     �?#       *                 ���2?.ݖv`p>=            p@$       '                 ��Dm? /y��C=             @%       &                 ����? � ��=              @������������������������       �                     �?������������������������       �       �             �?(       )                 ʊ�X? {�&��=             @������������������������       ��o�	��<             @������������������������       �                     �?+       .                 ��+p?ȿ���==�            �o@,       -                  �0��?�`\A=
             $@������������������������       ���q�4=	             "@������������������������       �       :             �?/       0                 `�݇?��]
��<=�            @n@������������������������       �Nh���!=             9@������������������������       ����Q�>=�             k@�t�b�F      h�hhK ��h��R�(KK1KK��h �B�  ��E���A>����V�V	�f��N����r�T� ����P�Bb�<��[�L�d�����ލB�O���d�><\e�VU�?���H��?��nVQe���vVU�K�pmUU��=��VU�?	Nz�{��9�f�����Յ�������UU忁uQ-VU��OK}UU��T4�i��?��UU�.�͆	N� ��^UU�`bv\UU�?t�W%A�`>��U��>�M��$��>���ZUU�j��VU�?����WU�?ps=�X>Z�C�VU�?ĂT�.#T>%w���~���w-�����c_sAVU�
67�VU�p�=n�d����UU�p�h}UU�?��:\>�����>\�I����?�&ɝVU�?N�.�
>T>b`N�w�´�� E�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K9h�hhK ��h��R�(KK9��h��Bx                          �@�F?}5r��J=�           �}@                        �HA?:��Sx�O=	             "@       
                 X�Oq?pg�L,N,=             @                        ��]?Hs�^�'#=             @                        � �5?�]�O�=              @������������������������       �                     �?������������������������       �                     �?       	                 ���`?������<              @������������������������       �                     �?������������������������       �                     �?                        �/5?0"$�~�<             @������������������������       � 2`�W��<              @������������������������       �                     �?                        l�*v?@���2=              @������������������������       �                     �?������������������������       �      0�             �?                         �ĵP?1���J=�           �|@                        ��g�?�I>�;=             (@                        ��IL?��o�;,=             @������������������������       �                     �?                        `�GM?(�ÿ���<              @������������������������       �                     �?������������������������       �      ȹ             �?                        0��?���3=	             "@������������������������       �                     �?                        �4Aa?��zHp4!=              @                         ��^�?x`�,���<             @������������������������       �Pt ���<             @������������������������       �      �9             �?                       ��ӉW?pI+Oǩ=             @������������������������       � ���$��<              @������������������������       ���o�D�<              @!       *                   �G�?*�h�J=�           0|@"       )                 �7~�?6�G{�L=<             N@#       &                 P]ڒ?
���?K=;            �M@$       %                 �/��?^���3Q="             A@������������������������       ���55W�F=             <@������������������������       �"ӆ^W=             @'       (                 0]�?.S�:�8=             9@������������������������       ����.�U=             @������������������������       ��$:�r*%=             6@������������������������       �      n�             �?+       2                  �P��?\�t�/AJ=�           px@,       /                  bB?)La�)E=G            �Q@-       .                 �f)??ٺ���GH=2             I@������������������������       ��
x�C=1            �H@������������������������       �      d:             �?0       1                  �0�?�gh�P� =             5@������������������������       �p6��WB"=             @������������������������       ����˕�=             .@3       6                   \��?-��K=@            t@4       5                ��G��?���+WP=	             "@������������������������       �h�k�J2=             @������������������������       ��G�4�D)=             @7       8                 �9a�?B`�J=7           ps@������������������������       ����8\T=a            @X@������������������������       ������C=�            �j@�t�bh�hhK ��h��R�(KK9KK��h �B�  j���e_O�w���\؎> I�'d'>@��{|q�>��� 4L���~UU�>�tUU�?  `�S�>�jײUU�?��I�UU�?�c�ީg��V?��UU��c�UU�   �0�>�Oo�VU�?
���VU�?��ں��T�@���񃐾-�m���u>ڔ��UU�?<j���t��[�xUU�k��hUU�mJfҗ� ßVU�^��� ��#-t9L^���b�UU�6JjUU�*03�m��puo�UU��VU�I����L����xw�y�ۭݡxnu�J��4�މ��(�<�ǿ@��VU����s>h dQVU�?�PU�W2���\�VU�<�ֲ�7���$�B�y>9c�;�>)�ǊQ:�?){vvWU�?x������s���UU���Q�UU�K��S�W�����z����BWVU�_�XGj�?Q�˟�L���!�j&�?�ڏ��Aÿ�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KQh�hhK ��h��R�(KKQ��h��B�                             �G�?��%U��O=�           �}@                        �7~�?~SO�#�K=@             P@                        P]ڒ?�Z.{J=?            �O@                        �/��?1r�"$O=&             C@                        �t?���$D=              @@                         a�U?�}��F=             2@������������������������       �
��Yj#=             @������������������������       �������I=             &@	       
                 ���}?�T A��7=             ,@������������������������       ����l�=             @������������������������       �^{Ō �8=              @                         M��?8pQ\uW=             @                        ���?  o�T�<              @������������������������       �                     �?������������������������       �      @:             �?                        �~1�?���x�q2=             @������������������������       �h�M%a=             @������������������������       �       �             �?                        0]�?��cI��==             9@                        �fA? !-�#!=             @                        Ї�?�kw]�:�<              @������������������������       �                     �?������������������������       �      (:             �?������������������������       �      8�             �?                        �ab�?�bJ580=             6@                        ��(�?�0A�u�=             @������������������������       ��G4�k%�<              @������������������������       ��V.�ީ�<              @                        0�~�?n�&�ߏ0=             2@������������������������       � �ng�N:=              @������������������������       ��1���#=             0@������������������������       �      n�             �?!       4                 ���;?L���P=�           �y@"       +                 PGT~?XZY[�S=4             J@#       *                 �g|?�4ח��Q=/            �G@$       '                 �U���B$tS��N=.             G@%       &                  .:q?ʹ�?�Z=             3@������������������������       � 2��'cY=             0@������������������������       �p�EA�<             @(       )                   E(�?-a�2�4=             ;@������������������������       �C�;5��F=             @������������������������       �"�uǻ#=             6@������������������������       �      l�             �?,       1                 @n��?��HTψ?=             @-       .                 �@�?��6-%r!=             @������������������������       �                     �?/       0                 �s6? � x�<              @������������������������       �                     �?������������������������       �       :             �?2       3                 H���?��Ne�=              @������������������������       �                     �?������������������������       �      �9             �?5       B                 @��t?��'��N=d           @v@6       =                 �jE?|�z��H=5            �J@7       :                 ��%f?X�/�bH=-            �F@8       9                 ��A?�M��W=
             $@������������������������       � �߷�г<              @������������������������       �����RU=              @;       <                 �x?�4'ln==#            �A@������������������������       ��Ó�)�2=             :@������������������������       �^:�F=	             "@>       A                 ����?�66��8=              @?       @                 F�e?\b��=             @������������������������       ��$(k�.�<             @������������������������       �L�0��<             @������������������������       �                     �?C       J                 ���`?שS4�qO=/           �r@D       G                 �m��?��y�C=             @E       F                  DA�? ��͏�"=             @������������������������       �X�����L<              @������������������������       � �ѡ�W�<              @H       I                 @�V?h��/{Y1=              @������������������������       �                     �?������������������������       �                     �?K       N                 ��b?�	��t7O=)           �r@L       M                 |m�S?0�:K6	<=             @������������������������       ����hI!=              @������������������������       �                     �?O       P                  �\�?$|C(N=&           `r@������������������������       ��U ���K=             (@������������������������       �����'�M=           �q@�t�bh�hhK ��h��R�(KKQKK��h �B�  u����B>AZ��~>i	�,�z>m��D~.�>��Nɺx>�b1����>��
�	�¿s��(��?��0�#h��V�UU�x"���7�?���clb�>  PF.u�>�c0VWU�?ahWU�?  x��<�>�_îUU�?L�gYVU�?����ve���՚[������M�8N;VU�h��VU���o|VU忐�x��h>  p0��>�2�UU�?e���UU�?9*��<=> �3VU�۹�B��?P���VU�?+n�ŭ�@��"�6z>J���� �>����>xT+��Δ>Le��J��?�|��UU忇@hU�JI>N�֞���?�K�DͿ:UK|WU�?�cs g�����C���7VU忲|j�PO��,�VU��]�VU忐�s�rYaO�UU��Y�pUU忡1 �f�X�ӷ�B�a��wc��:��6�LZ������VU�����ڿV.T���8�.gXt߿�����c�?E���w>�$�0ʼ�>���UU�?�~"�UU�?u�D@VU��H7���>�sI�Ě>�Z�(��>�">WUU忄��UU�?  ��X�>1��*VU�?���VU�?�(�_��?��9-6�4���XjVU�E��0WU�z����:!>?ʶ���2M�!�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KEh�hhK ��h��R�(KKE��h��B         *                 P�$�?��g:�&=�           �}@                        `���?�����"=�           �y@                        0<�?O!{���=<           �s@                        �R��?�X���=:           �s@                        0A��?B�%�q�=�            �o@                        �;�?v�1��`=�            `o@������������������������       ��t��`�=�            @o@������������������������       �      e�             �?	       
                 ���?x"}5�<=             @������������������������       �                     �?������������������������       �j�h`=              @                        PGu�?���	w-=<             N@                         `S��?`/�&!=*             E@������������������������       ���F3b�=&             C@������������������������       �ɽ�A�9=             @                          �x�?'��c��5=             2@������������������������       �<���L�=
             $@������������������������       ���{'�7=              @                        ��?��If��=              @������������������������       �                     �?������������������������       �                     �?       %                 ��]�? ���}�)=b            �X@                        pdJ�?����y&=^            �W@                          .p�?p��6S}'=)            �D@                         �1�?N�4z��<             @������������������������       ��Y(i��<             @������������������������       �                     �?                         �JV�?�8��&=#            �A@������������������������       �                     �?������������������������       ��BU�i ="             A@       "                 @� ?�ff��$#=5            �J@        !                 �8��?��r�I�6=              @������������������������       �45�r���<             @������������������������       �0�jo(%=              @#       $                 `�լ?�=-            �F@������������������������       ��V���)=              @������������������������       �QarŒ�=+            �E@&       '                 p���?Jq[kA�@=             @������������������������       �                     �?(       )                 ����?tZ!��s�<             @������������������������       ��?�-�!�<              @������������������������       �                     �?+       B                  �u��?�toːn9=:             M@,       9                 @8��?ĕ8���4=8             L@-       2                  �9��?4�\��qH=
             $@.       1                 �Vs�?�a$�(=�<             @/       0                  ��^�?Y,����<             @������������������������       �                     �?������������������������       ��F���$�<             @������������������������       �                     �?3       6                 K�ɀ?mĿ��K=             @4       5                 ���?@����=              @������������������������       �                     �?������������������������       �      0:             �?7       8                   ��?!�2�&=              @������������������������       �                     �?������������������������       �                     �?:       ;                 �=��?\�UW(=.             G@������������������������       �                     �?<       ?                 ���?�VR��&=-            �F@=       >                  ��?���4=             5@������������������������       �NHX7�	,=             3@������������������������       ��٦w�#=              @@       A                 �s�?&��Jb�=             8@������������������������       �]sҜ@ =             .@������������������������       �8�>'��<	             "@C       D                 ���?D{U��T=              @������������������������       �                     �?������������������������       �                     �?�t�bh�hhK ��h��R�(KKEKK��h �B(  Le�ZԢ:>�g� "���3u���R�"�Zѡ�O�I�;�_��@�vu_4�(��ř��HLU�UU�?   � �>CE+bVU�?��n�UU�?���E�s�q��qDP�C��[Gοp�Ԡ_��?Yr(�ŋ�EA̓�ѿQ��%����?�� ��V0�UU��֭-VU�[���q�j>�9@2�.e>�ծ� z>g�i��y�?�nUU忔�߸UU�]�q��q�>'�gVU�?0��˸�?4UT�1K5����
���p�9��vCq^VU�A�jB��c>D���UU�?̍z��?  h�b��>CF`�VU�?   �V�v>�zjUU�?����UU�?�Y�Q�p>��\w�h>�m9��e�>K�W�dQ�Z$i&��_��`vnUU���=_UU�ơxgUU�?  4Lp�>  ��m�>a��VU�?�iO�VU�?  �4�&�>
��UUU�?����UU�?
Ԅ	4/>]���UU�9�>�AJJ>H�YW
jp>��SK�?L�G0VU�?
i�3�f`���,?	俵��tUU�?  @��[�>���VUU�?Z���VU�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K?h�hhK ��h��R�(KK?��h��B�         >                  @���?��L��@=�           �}@                        @F��
�H�@=�           p}@                         �v�?a-���;B=�            �k@                        ��v�?��E�dD=y            @^@                        `�լ?%�	Dmh@=c            �X@                         �9�?Cq�A��8=             =@������������������������       �Y���=             :@������������������������       �T�T��=`=             @	       
                 0=T�?L��P��@=F            �Q@������������������������       �����M@=?            �O@������������������������       ����'U�1=             @                         ��?C�-���J=             6@                        `.��>_�#8=             @������������������������       �                     �?������������������������       �ƁdY)	=             @                         �g<�?����#J=             2@������������������������       �EM��a�)=             @������������������������       �0N�O@#K=             (@                        �g	�?�����==d             Y@                        L
�?�@M7
�(=             @                        �.�l?�f�
=              @������������������������       �                     �?������������������������       �      :             �?������������������������       �      "�             �?                        `���?I;h�R;=a            @X@                         ���?O�����H=!            �@@������������������������       ���H>D=             >@������������������������       ��h��_v=             @                        ��)�?�,��yt+=@             P@������������������������       �.�c�+=             &@������������������������       �<�i]�&=5            �J@        /                 �D�澙��͸>=�            @o@!       (                 �v��?�����E=Q            @T@"       %                   ��?��A�
D=<             N@#       $                 ���0?RG��=             @������������������������       �                     �?������������������������       �85���n
=             @&       '                 �c?�?�����B=5            �J@������������������������       �ӕ��NA=3            �I@������������������������       ��(Z_�,=              @)       ,                 p��?���d'7B=             5@*       +                  U��?4��-?K=	             "@������������������������       �.���<              @������������������������       �      0�             �?-       .                 �8d�?�u��ڥ)=             (@������������������������       ���Y��$=             @������������������������       ��s*Ti�<             @0       7                 �I�?��۷R7=�             e@1       4                  I�?��~H�K=&             C@2       3                  ��}?�~����4=$             B@������������������������       �t�,
J:=             0@������������������������       ���¸�#=             4@5       6                 �kC?:U˳m=              @������������������������       �                     �?������������������������       �                     �?8       ;                 ���?��co�?*=�            ``@9       :                  Ʉ?�VV_)kT=             @������������������������       �(+��A=              @������������������������       �                     �?<       =                 `I�?��"w/$=�             `@������������������������       ��t���:=             &@������������������������       �d��=u            @]@������������������������       �     $��             �?�t�bh�hhK ��h��R�(KK?KK��h �B�  N��Hdz2��47��98�-I���b��~�*�u��|�%�Z�����x>�����?�_ϘK�?��ܵs�c�K �ӿqT���?P�3I������~���.����VU�k�$�UU�?��J4?����(�F�ڿ�B��VU���
ʁX>UU&8]�>   �&�>;n{VU�?K�j-VU�?��#�UU�?|C:[p�6>r�(���{>k�:M~�?���nVU�?�_�bIuh����UU�:�v��&��q��n�U>e�:;z>�맜,�>=�����P�)VU忮mծUU�v���YW�>Sy�MN�?��6�VU�?ZR��?���3��j>L. �UU�(ܼWU�?�Y�����1���UU忍�P�UU��b�`�oR���Y�s>tQ�ԥ5>Z�0�m��?������  X~ѵ>�b��UU�?���kXU�?�!�RKg���ڱ�ߠ��̭�UU��^,WU����4�a����'���c?|ÿy`]5VU�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K[h�hhK ��h��R�(KK[��h��B�         4                 P�$�?��/ �sC=�           �}@       !                 ��{�?#�:�@2E=�           �y@                        @F�) 8W�D=�           Px@                         �v�?jQ�vF=�            �h@                        �G�?T�f{G=s            �\@                        -��?��#r8A=^            �W@������������������������       �W@
!z�@=]            @W@������������������������       �      y:             �?	       
                 `Fe�?Uoci�"U=             5@������������������������       ��c��Y�N=              @������������������������       �֐�S=             *@                        `I��?�h��C=S            �T@                        �$I�?���{��J=$             B@������������������������       �=N`{u7N=              @������������������������       �˛6D��E=             <@                        ���?-y+��'7=/            �G@������������������������       ���/l=�B=             4@������������������������       �g�Ī�=             ;@                        ��&�?4I<�.�B=�            �g@                         �9��?���{ F=q            @\@                        ��?
wKK1=             5@������������������������       �0�8i�=             @������������������������       ����� =             1@                          ��?�l����G=\             W@������������������������       �K+?4�Q="             A@������������������������       ������<=:             M@                        @3P�?�u���7=N            �S@                        ��?6����@=             @������������������������       � ���T�<              @������������������������       �    (4
�             �?                         �Β?��k�65=K            �R@������������������������       ��p��Z,=
             $@������������������������       �R���5=A            @P@"       +                 ���?���%G=             9@#       $                  '�?�Oìy�E=             1@������������������������       �                     �?%       (                 �c�}?P�����@=             0@&       '                  ���?L�7 |I=              @������������������������       �                     �?������������������������       �      �             �?)       *                 0�C�?2�z7=             ,@������������������������       �$��c@5=             (@������������������������       �l��U'��<              @,       /                 �_��?#`���%=              @-       .                    �?6��� =             @������������������������       �                     �?������������������������       � �)v�Z�<              @0       3                 `�r�?1Oh��=             @1       2                  `���?ֿ�U.��<             @������������������������       ����٥��<              @������������������������       �M�yAx�<              @������������������������       �                     �?5       F                 ��K�?�V=C�(=:             M@6       C                 ����?�sd4��%=             ;@7       <                 �{�?Ta墬�#=             6@8       9                4ƞ�?�II�u��<             @������������������������       �                     �?:       ;                 ��m?�J�}���<             @������������������������       �̧͡ʱ<              @������������������������       �                     �?=       @                 Ч�?��S��j!=             2@>       ?                 ���@?��7�	=             @������������������������       � ¡R�<              @������������������������       �`f����<              @A       B                  ���?�x���\!=             ,@������������������������       ��pm�X	=	             "@������������������������       ��<q��%=             @D       E                 `l_�?%:�'��<             @������������������������       ��ە���;             @������������������������       ��tnd�o�<              @G       N                 ��i�?����&=             ?@H       I                  �я�?��:#2=             @������������������������       �                     �?J       M                 ��?`v\K(*=             @K       L                 ���v? �w�[��<              @������������������������       �                     �?������������������������       �       �             �?������������������������       �     �:             �?O       V                 ���?�ط"+K=             ;@P       S                 ���?��}�55=             6@Q       R                 ��x�?c*�=	             "@������������������������       �Jp7M,��<              @������������������������       �      :             �?T       U                 �ݛ�?V�=���=             *@������������������������       �PA�=              @������������������������       ��
6�b<             @W       X                  PV��?=_�L�	=             @������������������������       �                     �?Y       Z                 �?��`0��<             @������������������������       ��B�8ت<              @������������������������       ��f�S��<              @�t�bh�hhK ��h��R�(KK[KK��h �B�  �ח��� ���mP;�A>�@�� 3�J��ni�Z>�E�ĵ�t>�ȼgC[>X$����?��NVU�G�����>�ڶʃ^�?��0
'��?9$r�sDi���N#1���n٭w�m�?�!|��ۿyk�*]�h>�2�w���?���יڿ����b��Z0'Hy�RoN�qv>�G��UU�b�q����?�!-0o���ٻr�ݿV~x�@*���C%R�+k>�=lv�>�e�\VU�?��sUUU�x�M�a>��R/࿷מE&�?Z�x��>:ի����>\h=�UU�t-M`H.�>  �f�ɫ>�0
WU�?�Un�UU�?}���>�/���?]����?6�O�}��u^h��r�=eUU�̆��UU�3g�=�(��;&8��i>���~UU�?�h�ZUU�+��UU忁Т2�t�e�D 6����1:��I�6g�0>�܅UU�?�!�}e�T��`UU�,ԇsUU忟�3m���
V=�M{�����UU忒iԷUU�K=�z_��dj㿻��u�|�UU忆��@	i>��UUU�˼�UU�?"�m�9uB��G�̽���XaUU�?��Um�g���m#�J��$V\VU応!3VU忨��jUU�,�Ԟu_>��oь;n>�<1]��U��Z�л俚��UU�?��D�Sa}>����L�?�^WUU�`?�)Ox�NɽUU忝�^��d����oUU�?pGZUU忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K+h�hhK ��h��R�(KK+��h��Bh	         *                  @���?e^f-=�           �}@                          p��?9!V�#�=�           p}@                        `r�t?l���=�           �z@                        � �J?�'�4�=S           0u@                         ��I?��)�k�=           �q@                        @F�b�勺�=           @q@������������������������       �S�J�$=�            `d@������������������������       �QL���=q            @\@	       
                 �i��?�"u��A.=             @������������������������       ��3��Q�<              @������������������������       ��'�� =              @                         �L?(�j��=;            �M@                        h��?���=ƫ=              @������������������������       �                     �?������������������������       �      �             �?                         �^��?�wK7<T=9            �L@������������������������       �a����=8             L@������������������������       �                     �?                        ��Cv?!��&��=Y            @V@������������������������       �                     �?                        `Q�?o��Z=X             V@                        ��L�?���X=7            �K@������������������������       ��$;�W=&             C@������������������������       ��y>��=             1@                        p��z?�Y��<!            �@@������������������������       �                     �?������������������������       ����WA�<              @@       )                 �2*�?̼7���=+            �E@       $                 P�bf?��K��=*             E@       !                 ����?kع��� =             6@                         ؠ�p?Q#�l+=
             $@������������������������       �+��|�<             @������������������������       ���N�	�<             @"       #                  @�9�?|L)�S�<             (@������������������������       ��E�;7��<             @������������������������       � ���L�<              @%       &                 ��r?<��u�=             4@������������������������       �                     �?'       (                �Ck�`?��ɸ��=             3@������������������������       �                     �?������������������������       ��=>祦�<             2@������������������������       �      B�             �?������������������������       �      �:             �?�t�bh�hhK ��h��R�(KK+KK��h �BX  7�dB�:>�B��>>��J�YV)>T�>H]0���CZ��<>�,�\(n3>e@���?��L�9ſ	t�]|�>3�{UU�$�e�UU�?c�����l���fkv���X,�VU忮 0�UU��7́�f� ��>��Ͽ%z��UU��ᆗT�^>7VU�?��y]�X>���vog>��}���?~xіUU�?[��D�GI�����UU���!Ӡ8��A�� j>T���wec>���9��;�,=��ջp���)oUU忒QբUU�UUUhd�e>��zUU�?C�bUU�?b�#Gv>�K4VU�?�h��lLm>�.;�UU�?�����?j�VU�?e��UU忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�Kkh�hhK ��h��R�(KKk��h��Bh         8                 �.��?��[SW/=�           �}@                           �?Q���2=#           0r@                        �F�f?�c��*=�            `e@                        ��??�k�6.=J            �R@                        P>�j?�+0H(�.="             A@                        �Ib?O�O�;@<=             *@������������������������       �����N =             &@������������������������       ��l��wx=              @	       
                 ��'|?�h94`?=             5@������������������������       ���9/�<	             "@������������������������       ��:�V��=             (@                          p��?�&�إ�*=(             D@                        ���L?�x|*�N(='            �C@������������������������       �xeJY֪&=             :@������������������������       ��xD�Ab"=             *@������������������������       �      S�             �?                        `|)�?M��&=a            @X@                          +Y�?X*ZԌ�2=(             D@                          .p�?�V���1="             A@������������������������       �-�xo�Z=             (@������������������������       �@�:�2�4=             6@                        �Ix�?��K���$=             @������������������������       �V�Z���<             @������������������������       ���l޹$�<             @                         �6�?�&�=9            �L@                         �x��?��&��"=             0@������������������������       �>���<             &@������������������������       �y�3Q,0=             @                        `��?�i?�3u=)            �D@������������������������       ���Xp	=
             $@������������������������       �*��IW��<             ?@        +                  �g<�?�߲��8=x             ^@!       &                 �{��?dT�Y!=)            �D@"       #                 ���>�,��i=#            �A@������������������������       �                     �?$       %                 @�4�>�fiC1="             A@������������������������       �                     �?������������������������       �N: ��=!            �@@'       (                  ����?��5��&)=             @������������������������       �                     �?)       *                  �3��?��!��=             @������������������������       �                     �?������������������������       � e���\�<             @,       3                 @��?�Z�N>=O            �S@-       0                  ���?L�r��N=             ?@.       /                 �j��?.}���XH=             =@������������������������       ��R1���3=             6@������������������������       ����0W=             @1       2                 p���?|��a,V=              @������������������������       �                     �?������������������������       �      ,�             �?4       5                 (�0v?�[���L=0             H@������������������������       �                     �?6       7                  /Ⱥ?��(� =/            �G@������������������������       � ���t��<              @������������������������       �Ϭ`��!=-            �F@9       T                 ��?�@����&=�            �f@:       E                  �g<�?�U�5w�4=F            �Q@;       @                 P���?���*=              @@<       ?                 h�37?J��j�5=             @=       >                 ��E�?����<              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?A       D                   \��?�v]��9"=             =@B       C                  �9��?24��� =             <@������������������������       �/��Xo==             9@������������������������       �XJ_f�2=             @������������������������       �      :             �?F       M                   �P�?�|� �9=&             C@G       J                 �/��?������P=             @H       I                    �?Fa���=             @������������������������       �                     �?������������������������       ����OO�=              @K       L                    �?��c�2=              @������������������������       �                     �?������������������������       �                     �?N       Q                 P���?���p�+=!            �@@O       P                   ��?��Ɖ�4=             @������������������������       �                     �?������������������������       ����*R�=             @R       S                 �W�!?(�A��%=             =@������������������������       �                     �?������������������������       ��q��!=             <@U       ^                 @8��?�N'�3==o            �[@V       W                 @�Dv?����R#=J            �R@������������������������       �                     �?X       [                 @�ե?��I@S=I            @R@Y       Z                 �&�?x�$��=             *@������������������������       �l%<d�=              @������������������������       ���ͫ���<             @\       ]                 �DT�?=Z����	=<             N@������������������������       �|O�5��)=              @������������������������       ��٭'�=:             M@_       d                 ��Q�?>W
�*�=%            �B@`       c                 ��F?$�.H-!=              @a       b                �٬Ӌ?��9ζ=             @������������������������       �                     �?������������������������       �@�����<             @������������������������       ���!�]��<             @e       h                 ��N�?��b��=             =@f       g                 �Nͼ?�3Y����<             *@������������������������       �c����<             (@������������������������       �      �             �?i       j                 ��ѽ?]��=             0@������������������������       �|�8��$=             @������������������������       �J�*�l�<             *@�t�bh�hhK ��h��R�(KKkKK��h �BX   E�9��S���Z���1��!>�L�Y�(m>�2X�9���O���%3ێx����mVU�$�G�q>��N�UU�?/)��#(�? ���<T|>yFF�:t>�{�q�?k��P�?3X�UU応/�"�Hd�}�ڵ54v�y�?Fc!��,�ܒ��?JA�࿷[:�d�>:�ہUU�_�UU�?x�ۙq�:�M(h��k>gb+ЎLӿ���C4�?�ʭ�_�ZZ@�UU��$L@r�?���q�W2i�Z>��#�P�&��9$�UU�?��>xP���a�UU�e�*�a����;Μ�>V�~!VU�?�u-~r}>����UU忻�c�UU�?��\�&i}��zBIp��IL��9߅��d���ǿU��VU��Ǹ��鮾���gWU��&+�UU��XޙXg��W�!VU忡����Ra�� ��UU�?X������̐��Z>���u>L���O">�w�H]��0.#���|�f�`qUU�d�\�UU忹]NVU�GCN �b>����i>v/=�d��?��pD�?��a�UU�j�q�-�>�Z���5�>�g�:|v>f���UU�?'�#�S즿  �ư>���^VU�?�!�WU�?�$�y>  (�쵖>�pC`VU�?�Mf�UU�?�́I��p>���UU�5�׳���?�sM_�B�>�L�'_�����UU�?�P8�f�a�,�P�T��̎#��ܿ ��UU�w�g�+O��p[k?�?(7N�x�ӿ\lv��`>��\i��>  ���>�VU�??&��UU�?�9]UU忹ד�νM����b�p�xgUU�E�y�UU�A�¹:�^>>Rqt�x�?Z����ϑ?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KWh�hhK ��h��R�(KKW��h��B         "                 ��cn?r$Y�2=�           �}@                        @淨?~�1�f:=C            �P@                         խ�?�X����5=;            �M@                        ��?0���52=8             L@                        P.�?V7�i�:=             8@                         m�a?}���m+=             5@������������������������       ���-;³!=             0@������������������������       �����Q�!=             @	       
                 ��	<?�3�}8=             @������������������������       � híE�<              @������������������������       �      :             �?                        �x�?�LEw�Z$=              @@                        ����?���� !=             >@������������������������       �q��k
=             9@������������������������       �	�e˧#4=             @                        �da?`��9�<              @������������������������       �                     �?������������������������       �                     �?                        t��?T]JT��4=             @������������������������       �                     �?                         ��?@t�?�<              @������������������������       �                     �?������������������������       �       :             �?       !                 ��p�?|���3(I=              @                        pz�o?qe�p0=             @                        ���`?7�-#3�
=             @                        (;Ja?�Yͷ��<             @������������������������       ��7�
1�<              @������������������������       �                     �?������������������������       � ���9|�<              @                            �?l�ib 5=              @������������������������       �                     �?������������������������       �                     �?������������������������       �      0�             �?#       :                  �kI?�l�ˁ1=�           Py@$       1                 �x?�n�^�*=:             M@%       ,                 @*tC?��Ȝ9i"=0             H@&       )                 0��> u���=*             E@'       (                   ��?9hOZ�=              @������������������������       �~X{�U�<             @������������������������       ���*�~#=              @*       +                  `���?����<="             A@������������������������       �E�v=�=             @������������������������       �����.C=             ?@-       .                 �g�G?&�<t:�+=             @������������������������       �                     �?/       0                 P�n?d���`=             @������������������������       ��J���<             @������������������������       �      �9             �?2       5                 `�@|?�g]	;=
             $@3       4                  �Q�?�4�6n�=              @������������������������       �                     �?������������������������       �      :             �?6       9                 �NN�?���7��=              @7       8                 8���?(r.��Z=             @������������������������       �L|�ߩ��<             @������������������������       �                     �?������������������������       �                     �?;       H                 �SpR?i���>�1=[           �u@<       C                 ����?�@nxC=             5@=       @                 �=l�?r:���D=             0@>       ?                 �u)�>����$=             ,@������������������������       ��];���=             @������������������������       �<��X%=	             "@A       B                 ��Dm?����^=              @������������������������       �                     �?������������������������       �      @:             �?D       E                  A��>�ԫ��d=             @������������������������       �                     �?F       G                  ����?\0X�9�<             @������������������������       �                     �?������������������������       ���C�
�<             @I       P                 �\ͥ?*Yս4i0=F           `t@J       M                 hU�<?����v4=              @K       L                  ���? �1:k�=             @������������������������       �                     �?������������������������       � *��<              @N       O                 h�b?�D�a*�<             @������������������������       ��*����<              @������������������������       �KhC�X�<             @Q       T                 `��?���3t&0=>           �s@R       S                 �%�?��f�ql>=             &@������������������������       �                     �?������������������������       �i�'L(=
             $@U       V                 P�Y�?�o�Å�.=3           0s@������������������������       ��2�K=             1@������������������������       �^j<�h�)="            r@�t�bh�hhK ��h��R�(KKWKK��h �B�  ��:�J>.��!�g>"��3�T>�8^�x@g>�ĕ8�.�>�-	��g>�%���¿@Ԗ�UU�?UU5���>c)k�VU�?/���UU�?̨q|roO��צ_�c��A��?��'���  �َ�>��UU�?���UU�?e#i(�����yVU�~c��,�����UU�'��UU�8��]���>�`��m�x>�`����J��T��m'q>9�kF��?"*��UU�?{�UU�  PV��>�euqUU�?*G5VU�?���VU�?��]A�6��O��q�-F�H�y�׌'T��K7
ǟ9�{l�rUU�,W �?3��T����D֙��?zB��UU�ݐ�6x>��VU�?���o�)>�K�>(��?���UU�
�n's>  ��ʙ�>��SVU�?N��VU�?t.�r$rq�W�8[�W����?��'�UU��w�UU忮�Sb��4>u�@�>0���6�>�+ �u}>��KI�@���5�UU�?  P����>6���UU�?��HsWU�?S�C���W"�UU���o�m�� (\UU�?��sUU���G��)�jU�>������������?VU忾�y�UU��3���g>�<Q�UU�?���^UU�Y�d��d>6e�X�x�>��~�VU�?�oSQD�?���'�5����{+��?�n������t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KEh�hhK ��h��R�(KKE��h��B         :                 �)�?�`��L�=�           �}@       !                 0vb�?;cm�v=�           �|@                        0��?%}��=�             o@                        ���?艁[4�<�            `a@                        pb��?��Z~z��<�            �`@                        ��m�?irVT�<w            �]@������������������������       �8��陟<u            @]@������������������������       �|�6Q5U�<              @	       
                 k�?��x�d�<             .@������������������������       �                     �?������������������������       �ٱ���<             ,@                           �?��	���'=             @                        �_��?x;̐~=              @������������������������       �                     �?������������������������       �      �             �?                        `l,�?O�j:�{�<             @������������������������       �                     �?������������������������       �  �� <              @                        �\ͥ?5����w!=n            �[@                        (�e8?��[�Å4=             @                         ����?𠏶�3=              @������������������������       �                     �?������������������������       �      �             �?                        n�
Q?�##y{q=             @������������������������       �p�ߝW�<             @������������������������       �� }�Ƽ�<              @                        ��Ҧ?�~�\x=g            �Y@                        0Du�?��b!=M            @S@������������������������       ����o=@             P@������������������������       ��W��R43=             *@                         `Fe�?}FK(�=             :@������������������������       �Ǎ�ZX�=             8@������������������������       �D�L��=              @"       /                 �7��?nCe}8:=�            @j@#       *                  �8�?4����:=�            `e@$       '                 `�0z?�i� ј=�            �d@%       &                 p� �?mE��=�            �a@������������������������       �O���F =            �_@������������������������       �3�4=             *@(       )                 @u�?���a�<             :@������������������������       �8�_�&��<             @������������������������       �����C�<             7@+       .                 Pα�?�ʇ��*=             @,       -                 d�?�?�¶��=              @������������������������       �                     �?������������������������       �       �             �?������������������������       �����f�<             @0       3                 8~U�?>��r��<'            �C@1       2                 x�b�?@gƇv=             @������������������������       �h]X�Ԑ�<              @������������������������       �                     �?4       7                 @��?�;ZQ��<$             B@5       6                 �9��?X�����<             ,@������������������������       �H��c��<             @������������������������       �g�~�N<�<	             "@8       9                 p[͔?���:b1�<             6@������������������������       ����Ƀg�<	             "@������������������������       ��l ��I�<             *@;       >                 4 �?,?,<:=             *@<       =                  >��? �uL��<              @������������������������       �                     �?������������������������       �                     �??       D                 ��?lw�&��<             &@@       C                 @���?��~R��<             @A       B                 ����?�����3�<             @������������������������       ����D�<              @������������������������       �                     �?������������������������       �j-(���<              @������������������������       ��))`�|<             @�t�bh�hhK ��h��R�(KKEKK��h �B(  JpC�\2>i���d#>��-d>G>yqB H�4��0���F���ط�:��<�_J��E��UU念��/hi���%�UU�5pIQ;���w���>  P�gq�>#"j�UU�?��	VU�?+M7W��#>@��nUU�R�\cUU�?��5l`>h�?ʄ>  ��ja�>��KVU�?��!�UU�?M�b�4a#�/�=˘�`��UU�?��� �W>
m͒[�d>e��[��?O�}��?��#+/X[���D�ڿ3�UU�?LՐ��@��.ii��O�x6�K�G��e����U���`��ɿc��^{��vb'�ed>1Y��UU�?Z��eUU�?k#JZ�m��F��Lݘ��s�UU�=��VU��t^]UU�?0�ݮW>UU�M��>� bUU�?��`�UU�? QJM��L>�m[ѫ�a>���wUU�?-�\UU�?�4kX�>J�bUU�?,����׿�R�R�s>  px��>"��UU�?&��UU�?\u�3xY>�����k>����ut>o��kUU�?�zUU�?H�]UU�?q��^
y�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K3h�hhK ��h��R�(KK3��h��B(                          h�[�>LЁ]=�           �}@������������������������       �                     �?                        �`>R?:z��=�           p}@                        ��IL?
%�=             6@                        ���J?J�:�=             (@       	                 �@�F?N��R��<             &@                        @{d??���.?�<              @������������������������       �W����(�<             @������������������������       ��O�*.�<             @
                        X�D�?��k"��<             @������������������������       �                     �?������������������������       �h�c_�K�<              @������������������������       �                     �?                        ��f?�h?�K)=
             $@                         ����?�+ȩ�<	             "@                        �U�?
���d�<             @������������������������       ��k��S�<             @������������������������       �      �             �?������������������������       �X5�&[�<             @������������������������       �       �             �?       $                 P�}A?eMw��=�           |@                        �&�?tՋg�%=�            �o@                        `Zf~?f���'=�            �g@                        ����?�҇��=�             b@������������������������       ���_��=Y            @V@������������������������       ��j�s\q=8             L@                        �X\�?(����.=+            �E@������������������������       ��d�ǟ=*             E@������������������������       �     �2�             �?       !                 �Y&�?x�q4==@             P@                         �=�?ķt�v.=              @������������������������       �                     �?������������������������       �      �             �?"       #                 @��8?λ�7�j=>             O@������������������������       �/6�6�<<             N@������������������������       �XN,�Ee=              @%       ,                 P�$�?��y>l=�            �h@&       )                 @�q?<;��<g            �Y@'       (                 (��?�2M
N=:             M@������������������������       ��� cT�=+            �E@������������������������       ��Ҫ�Q=             .@*       +                 �ގt?���:�<-            �F@������������������������       �                     �?������������������������       ���;-�<,             F@-       0                 ��?k!1�fn=^            �W@.       /                  ��?,�ֽ��%=             3@������������������������       �F�d�S0=	             "@������������������������       �UI� �<
             $@1       2                 � v�?��5~��<K            �R@������������������������       �,�n���<1            �H@������������������������       ����#7��<             :@�t�bh�hhK ��h��R�(KK3KK��h �B�  ��4' ��e��UU�?f}&	�#����q�h��hFS�y>�a�=�<W���j� .>^�K���࿞�yUU�?3%����w��gΌUU�&�6kUU�(�g�UU�?"9���{�� ,� t��g��9O�Q��{UU��:��UU�s@�^UU��
q�UU�(t����w!�cB>Ȅ
`rZR>':�k��8>�_���U�?�����˿�	#:�m>�|��:��?�>��UU�)4�R�Q����5[���)%VU��ԣ~UU���k�8�.��ɿ(U&�UU�?a�'�;H�R�iS��_�v&i�rk���@�Կ"��UU������#�9�InUU�?�#jUU�K��I�>C>����w>�
L���?>��Q{��?rI�F`H�1�����Q����T�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KSh�hhK ��h��R�(KKS��h��B(         *                 P�$�?|����=�           �}@       !                 0���?�	zs��=�           �y@                        ��?�����=�           �y@                        `���?�1�xɜ=           q@                        �kd1?�T
�[=�             n@                        `Zf~?���c�==�             a@������������������������       ��ڎ(�=u            @]@������������������������       ���0�P�<             4@	       
                 ��?n$�oܳ=h             Z@������������������������       ������=T             U@������������������������       �$��_�#=             4@                         �^�?LV#7�N=              @@                         �g<�?���D�+=
             $@������������������������       �����ֶ<              @������������������������       �Q���$�<              @                       ���q?�Ὀ��=             6@������������������������       �g���6� =              @������������������������       ��G���<             ,@                        @�ե?���
=�            �`@                        'm�?��+Z�%=             4@                         v_�?������=             .@������������������������       �Q�/\=
             $@������������������������       ��0׬� =             @                        ����?��A�G=             @������������������������       �                     �?������������������������       �h���y =             @                         ���?���=s            �\@                        �<�?h+�zT=	             "@������������������������       ��.0�t
=             @������������������������       ��iJ��<             @                         �<m�?�^�F�=j            �Z@������������������������       �vrǔ�u=             9@������������������������       �_ɤ��=Q            @T@"       '                 �V��?�e�V��=             @#       $                    �? ���	=             @������������������������       �                     �?%       &                 �F��? � ���<              @������������������������       �                     �?������������������������       �      �9             �?(       )                 `�r�?�x�f�z�<             @������������������������       ��!#�b�r<              @������������������������       �                     �?+       @                 �Y�?~�y��<:             M@,       1                 \��X?�Ӌt��=             ?@-       .                ��>T_?�,�{��<             @������������������������       �                     �?/       0                  `%+�?����oӷ<             @������������������������       �                     �?������������������������       ���d�B9z<              @2       9                 P�s�? >�u��<             ;@3       6                 �(�?���~���<
             $@4       5                  �a�?���0��<             @������������������������       �Ǫ����<              @������������������������       �h�]�ο�<              @7       8                  �Z�?�zp��<             @������������������������       �                     �?������������������������       ���Ո���<             @:       =                 p���?}aЁ��<             1@;       <                 nn?ℋ��<             &@������������������������       �
�픉�<             @������������������������       �,b7�L�l<             @>       ?                 P'��?~�+���<             @������������������������       �                     �?������������������������       ���x��<             @A       J                 ��K�?]qe9:�<             ;@B       G                 ��G�?�����<
             $@C       F                 �H��?����<             @D       E                 �=��?"A}c�<�<             @������������������������       ��(��5�<             @������������������������       ����fDd<              @������������������������       �      й             �?H       I                 p4N�?�w5QU"�<             @������������������������       �                     �?������������������������       �b�bPQQ<             @K       P                 �s�?O>&���<             1@L       M                  `���?��m���<              @������������������������       �Ƈ�&�<             @N       O                 ��s�?@+��W�<             @������������������������       � �	?[�<              @������������������������       �                     �?Q       R                 �r��?b��Q��<	             "@������������������������       ��$g���Z<              @������������������������       �                     �?�t�bh�hhK ��h��R�(KKSKK��h �B�  �a�@T�=�!5�	1>F	���#>������:�u����R>�~�,�Q�����Á���eZS���j��l�[>B��@�?�2k8��?dx��"q�^�x�`>�;ޜUU�?�x�56f��`�U�ΐ|�\$��UU忕�aq�係s`-U>^�����>,�A���j>u�E���?����}J޿��L�,�>)(�0VU�?6���UU�?_v^i+>��}ٮ�}���(�ːɿU��UU忡���H>�Qg���?zWCSA��_�K��>UUu��Đ>E��UU�?  �20��>��#�UU�?K�7�UU�?h����_S�>�FXUU���)eUU忴Cҋ\���N�Vi�0%�8Q6i>�Zq�UU�?��u~R>Zg]dUU�?ZȃQ�?�M��ip�}�b�r��(��ƺp�ʵ�yUU��`UU��*�*օ��X��UU�
�~�UU忮_4|�Z�Q��n��FR�UU忯�PXUU�b �y
a>�w΁UU�?�F>��?	�0-� �MXPLL�[���1N$j�gZ8��M`���3hUU忨��WUU�m���UU志3�W��B>0{�cUU�?��VUU��8BYO�I>�f���eb>{�����?UUՈ�v>$*nUU�?��e�UU�?���-�@��"WUU忶��gUU忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K-h�hhK ��h��R�(KK-��h��B�	         *                 ���?"Uk�F�<�           �}@                        0���?z�-��<�           `}@                        ���?㽓 ،�<Q           u@                        P!d�?�PN��%�<M           �t@                        ��y�?�F{��e�<>           �s@                        P�,�?�39�T�<�            �m@������������������������       ��n�uQ�<�            �m@������������������������       �     @7:             �?	       
                  �?y�!'5�=Q            @T@������������������������       �                     �?������������������������       ��<l���=P             T@                         `S��?.��z��=             .@                        ��H�?4ԁ>O��<             ,@������������������������       ��5&�c�<             *@������������������������       �      �             �?������������������������       �      �9             �?                         �E�?e�w���=             @                        �m��?�m[�q��<             @������������������������       �                     �?                         ��?��]�n�<              @������������������������       �                     �?������������������������       �      ��             �?������������������������       �                     �?                        @K�?�)<��<�            �`@                         ���?(� ���<              @������������������������       �                     �?������������������������       �      ع             �?       #                 P[)�?|����+�<�            ``@                         |�L?��S�} =             0@                         �P�?�m~��=             @������������������������       �                     �?������������������������       �,�no8�<             @!       "                 ����?�.;[��<
             $@������������������������       ������~�<	             "@������������������������       �      �9             �?$       '                  �~��?o`4�W��<s            �\@%       &                 �$I�?�%:�ml�<             <@������������������������       �                     �?������������������������       �u�ݔX�<             ;@(       )                 `��?����7P�<W            �U@������������������������       ����ND�
=              @������������������������       �Q����<U            @U@+       ,                 J�$�?�ut �=              @������������������������       �                     �?������������������������       �      �9             �?�t�bh�hhK ��h��R�(KK-KK��h �Bh  �z�>�>V}�)?�>�ޣ,1%�N�\Wy��@

�}>�@IU~0�H丩�ſ}�АUU�?�^|BS>eE"�UU�?͜B��@�?�gdZsj���u¸Er��`| 忩�%�UU��MR�UU�?y���4���B��cqs�&��UU������Z�^VUU忶��fUU�����UU��d�W1|F>  ��O*�>�UU�?�S�~UU�?������@>�*���f>��*��}>M���UU�?�M{{UU�?"�wrc�>!���`C�j�kUU�?<�
��*>�@w��qT�+�9�UU�B����ѿ�c��PF>��)��߿'K)]�:�?  @�(sz>�YܛUU�?�VUUU�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K-h�hhK ��h��R�(KK-��h��B�	         ,                  @���?�<^c�1=�           �}@                        �94W?⟹���=�           p}@                        ��bV?bQ1��=[            �V@                        �U�����͊و=Z            �V@                         e	a?ݴ���~=$             B@                        �$?Z?��d�=             0@������������������������       �T�v(/�=             *@������������������������       ����)���<             @	       
                 T�@?~<�顟=             4@������������������������       ���ef��<             @������������������������       �آ��D}	=             .@                        P^N<?kX�u��<6             K@                        �
OW?m�!Ї��<#            �A@������������������������       �܃��2I�<              @������������������������       ���a�A��<!            �@@                        P^�?�p֒�<             3@������������������������       ��L�v>�<
             $@������������������������       �#�{n�U�<	             "@������������������������       �      ":             �?       #                 ���u? ��I5�=|           �w@                         �_�?7$u��H=7            �K@                        ��_i?���H�=             ;@                        �p�?�u2ۼ�<             0@������������������������       ����m�<             .@������������������������       �      �9             �?                         ��i?V��ۂ��<             &@������������������������       �                     �?������������������������       ���<�l�<
             $@                          ;��?rȲ_�d=             <@                         `���?g��W =             ,@������������������������       �d�䡝�=              @������������������������       ���hG�(=             @!       "                 �&oh?bq�p�&�<             ,@������������������������       � �!z犿<              @������������������������       �mN�B���<             (@$       %                 0Vtv?����T)�<E           Pt@������������������������       �                     �?&       )                  �|?[��5�<D           @t@'       (                 h�2�?i�@@��=
             $@������������������������       �*��TL�<	             "@������������������������       �                     �?*       +                 �$�|?��TZ�N�<:           �s@������������������������       �                     �?������������������������       �7�5q��<9           �s@������������������������       �     �f�             �?�t�bh�hhK ��h��R�(KK-KK��h �Bh  6[�y	 ��t���$�\}��\T�^E��WQ��(ݭ�g��?��sT>|-���6ؿ���UU�?�_�R�y��A2�UU忛_%�	=��nd�X�&>o\>�?{`>�n��E�ZnUU�?\��OSj��Ű�.?俻��p_�?.���UU忢�~���>�C0.�b>�s�Ա�Q�oL��]>Б��3�?��UU忡��J�u���%�UU�<1X�UU��B~��v>Ւ*:\�>+9G�UU�?�=>���?���RU>2��UU�?qYTG��?��/?YT1�Έ��UU�^����(�Fg��Jq����	z�ݿ="�UU��~3�����0�UU�?���f����rG�UU�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KYh�hhK ��h��R�(KKY��h��Bx         "                 �94W?[��P�"	=�           �}@       !                 ��bV?��$E@;=[            �V@                        �U���T�\V�=Z            �V@                         e	a?�;�Jsu=$             B@                        �$?Z?l���E�=             0@                        �R$X?��$d�=             *@������������������������       �]�q����<             (@������������������������       �       :             �?	       
                 P��[?`"f0r��<             @������������������������       �                     �?������������������������       � �$����<              @                        �$܀?.���=             4@                        J%�?��:�=             0@������������������������       �d��gK=             .@������������������������       �     �)�             �?                        hpr�?d��.��<             @������������������������       �`�&��w�<             @������������������������       �      ��             �?                        P^N<?��R[,��<6             K@                        �
OW?Z�K��<#            �A@                           �?�CY���<              @������������������������       �                     �?������������������������       �      ��             �?                         P���?����-�<!            �@@������������������������       �                     �?������������������������       ����{T�<              @@                        ��V�?"ḻ"�<             3@                        p��W?�~�t���<	             "@������������������������       �                     �?������������������������       �$D	����<              @                          @(B�?vJ�2?�<
             $@������������������������       �8_�-��<             @������������������������       ���g��<             @������������������������       �      A:             �?#       <                 �pur?�fz��=}           �w@$       1                  �_�?��9~8=-            �F@%       ,                 0vb�?�X�7�:=             9@&       )                 P$�?'���^�<             6@'       (                 �2i?AT4
��<             3@������������������������       �s�{�n�<             *@������������������������       �Џ�X�
=             @*       +                 ���g?��H�-�<             @������������������������       �                     �?������������������������       � �c|*��<              @-       .                 �i?ȸ�!M�<             @������������������������       �                     �?/       0                 H^[�?x3�j�<              @������������������������       �                     �?������������������������       �                     �?2       7                 @��p?q'Nr�6=             4@3       4                 P��W?ӣ�F'd�<             1@������������������������       �                     �?5       6                 wr?$n
s���<             0@������������������������       �pVzs{s�<             @������������������������       �
Y����<             &@8       9                 \F�M?t%�'Ҿ=             @������������������������       �                     �?:       ;                  P�"�? �r:���<              @������������������������       �                     �?������������������������       �       :             �?=       J                 ��{s?�-��=P            u@>       E                 `��?�'�A;�<             9@?       B                 �m��?,�I,�. =             1@@       A                 0{l?&/���<             *@������������������������       ���_a�<
             $@������������������������       �P��F�<             @C       D                 pmgw?����bi�<             @������������������������       �                     �?������������������������       � �'C��<             @F       G                 �2N�?�|Ei:�<              @������������������������       ��{�΀<             @H       I                 ��8�?�
$L�<             @������������������������       ���!�T��<             @������������������������       �      �9             �?K       R                 �?���/�=7           ps@L       O                 Pc�?�=�;F�=             @M       N                 ��3G?[�_p�<             @������������������������       ���D��Ġ<              @������������������������       ���cGK�<              @P       Q                  ����? H�,?�<             @������������������������       � &�l�P�<              @������������������������       �       �             �?S       V                 �<�?�Z2�U&=0            s@T       U                 ��*?����	=+            �E@������������������������       ��
+=�=             :@������������������������       �sQ���=             1@W       X                 0�Z�?��Su9�<           Pp@������������������������       �I�
gZ�=>             O@������������������������       ��;�2	�<�            �h@�t�b��A      h�hhK ��h��R�(KKYKK��h �B�  �XHQ4�>�3��|�S>?�F��P>t�N���j>�K���S�>	rԸ�g>�!Vg��?��E�UU�?>�Lm`����zh�UU��w�UU��4@+|>#�,��с>Rz"���?y�rUU忍q%vv;�ݩj]UU�baUU�?b�g�:@��f&`�)���%Tk>��SUU�?{��ZUU�MRg���b�
Ph�UU�JY�kUU��\�	8b>Y$@�y>��M^UU�ݝ�UU�?~V"��V�Y,jUU�?M �mUU�ζUU�?���]i/��[w {h��k�K�AD�Q�.x��Y�x�̭P�D����?��������?X�(8�bڕgUU�`̊UU快����2z>}�z�UU�?  @g�]p>m^�_UU�?4@�vUU�?�.+5`x����	5bp�éD�UU忻Tl�@�i����UU�BVxʤԿ[?�]�j���+�aUU応!������UU�����UU忨6Q�3!>�d�
k>z	����t>f�C�G�g>�3�r��?�Mw�UU�?   �I��>G��gUU�? �UU�?�m��Bk7��݉eUU�?����c�J fUU�F">WUU�?��v��B �~����y�����?J�}2�cUU�0{\UU�?h��©��/,�UU�jv.�UU快��V��=^`�rd>F��Q�|��#>��Ƅ�?�����9���F�(�ҿ�K)�/�?�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K-h�hhK ��h��R�(KK-��h��B�	         ,                  @���?K��_��<�           �}@                        ��K�?���C�r�<�           p}@                        ��_�?���}t��<�             e@       	                 �j"�?`X�����<�            �d@                        P^��?���[� �<Y            @V@������������������������       �������x<J            �R@                        @F�� t�;1�<             .@������������������������       ������<             @������������������������       �wB��,�<	             "@
                        �}��?B�-�1�<M            @S@������������������������       �                     �?                         ���?X���<L             S@������������������������       �;�lX���<             =@������������������������       �Y�X}`��</            �G@                        `?fbz��� =             @                         h��?@d�ht2�<              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �9             �?       #                  ���?���D<�<.           �r@                        ��g?Mp3�i�<�            �n@                        �C�?���:�<�             h@                          Y��?�U^����<�             e@������������������������       ���'�K��<�            �c@������������������������       �~��9l�<             &@                        �vQ?@qԇ��<             9@������������������������       �6)�J��<             .@������������������������       ��>�.���<
             $@                         p�m?e8Ȫ�u�<4             J@                        P���?��`��M�<             @������������������������       �                     �?������������������������       �@��<G��<              @!       "                 @���?x�DI��<1            �H@������������������������       �~qτt�<             6@������������������������       �zs&�9��<             ;@$       %                 ��?$oD����<9            �L@������������������������       �                     �?&       )                 ��Q�?�;y�j��<8             L@'       (                 p��?���a��<             =@������������������������       �v)�Ab�<             1@������������������������       �\�X�z�<             (@*       +                  �w�?]j��R��<             ;@������������������������       �  ����<              @������������������������       �&�gjȝ<             9@������������������������       �     @L:             �?�t�bh�hhK ��h��R�(KK-KK��h �Bh  ��jY�>&0M��>�U�I��G>��^�B>�����2�.	��ٿ�̒���V��G[yUU�㕾��x��CBq�c�X>X��UU�?�QAMT>�b��vr��9v�U]o�?UUU<4a�>   ��>�>�y�UU�?w�/�UU�?�M�aUU�?��8TZ�.�2�r�=������xG��*A*�?�*��Oֿ(X�L�?��R?��b�t�hr�2�)�7��?�~��@>UUUw+�>���pUU�?����UU�?�UB�g��\eT�95�?�'͋��ѿ�"���vG>s���UU�?����cB>w:/U>-�fiUU�?RH&�_�?Z_��,�0ҌwUU�2���`C�?F��UU忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KAh�hhK ��h��R�(KKA��h��B8                          ��IL?�����A�<�           �}@                        ���J?��

��<             *@       
                 ���k?�Zi�v�<             (@       	                 hì+?.��k�<
             $@                        �PAC?vqo�\��<             @                           �?C�b ���<             @������������������������       �Z:�8�f�<              @������������������������       �x�!e�Ѓ<              @������������������������       �                     �?������������������������       �tJ̓��<             @������������������������       �  `4��x<              @������������������������       �                     �?       ,                 @�C�?Z�+Ix��<�           �|@                         �~��?:Ǌ��=�<H           �t@                         �ڦ?{B#�K�<{            �^@                        ���G?�TEGF�<O            �S@                         K�?� �;*�<=            �N@������������������������       �]�"��<.             G@������������������������       � ����m=             .@                         �9��?�m�d���<             2@������������������������       ��/��g�<             ,@������������������������       �l�Ѝ�#�<             @                         m��?ZX�]���<,             F@                        ��7c?|z�ם�<             3@������������������������       �P��:��<             @������������������������       �fn����<             0@                        �>}?�fج�<             9@������������������������       ��N���<             @������������������������       �����?�<             6@       %                   �P�?�{۱�<�            �i@       "                 �m��?�����O=
             $@        !                 P�Dv?#4O/+�<             @������������������������       ��&F�!�<             @������������������������       ���+�U��<             @#       $                 p]�?6���=             @������������������������       �P����<              @������������������������       �    ���9             �?&       )                 �-�?[�-�j�<�            `h@'       (                 �<�?�����<o            �[@������������������������       �T�΁�&�<]            @W@������������������������       �M���y�<             2@*       +                 ���?�jܫj�<T             U@������������������������       �                     �?������������������������       �%��"���<S            �T@-       4                 @�Dv?�����W�<�            ``@.       1                 ��t?�����k�<              @/       0                 .�X?}�Iva/�<             @������������������������       �,Y4��<              @������������������������       ��zT�8�<             @2       3                 8���?��F0�=�<              @������������������������       �                     �?������������������������       �                     �?5       :                 `�0z?Wb�����<{            �^@6       7                 ����?y��p�=             @������������������������       � ���Nl�<              @8       9                 �=�e?/ŕ<             @������������������������       �                     �?������������������������       ����7<             @;       >                 ����?f�/��C�<u            @]@<       =                 �p�?�n_�X�=             @������������������������       �N� �E��<             @������������������������       �                     �??       @                  5�?�K~Z#�<n            �[@������������������������       �f]��~�<(             D@������������������������       ���а�<F            �Q@�t�bh�hhK ��h��R�(KKAKK��h �B  _ޔ)���pr�� a>���y�+P>reXs>b'`�V>�����>�n�^UU�5��\UU�?�ϛxUU�?�f�_UU�9��sUU�?O���UU�?�����X"�t}�%5��H�;6K���L�pu.�2rU-d�>>��]OC��1ͶP$��?a=Y��we�A鵋0�|Di�UU忆1$��2_����Dp�i;�з�?���UU�L���5����F���?c���pۿcM�#��񽍡7���k>
��`�G>BR|�U�?K2�kUU忪Vo����>�H}�UU�?y�VUU�B,��)� ��->��LW���!��b�?`%_�3"H��$��UU�]�oUDYῗ&��î4>Jdd6rk>�m�^};>W��]UU忲�*�8�?  ��b�>u3��UU�?M��UU�?�X&��>�A�0�@s���_�UU��� E��1�bUU�=C1VUU���4<�7>���f��l>��ԨX_�?s���UU�?��� �h%>
P��¢�?/Z;��ǿ�t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�KIh�hhK ��h��R�(KKI��h��B�         ,                 P�$�?��M��<�           �}@                         �/�?^�g���<�           �y@       
                 ��IL?@�؃�0�<�           �x@       	                 ���J?��މ��<             (@                        ���k?�gea$��<             &@                       �&�Ye?�罂��<	             "@������������������������       �%����<             @������������������������       ��B`x�[�<             @������������������������       � �s�|�x<              @������������������������       �                     �?                         �~��?T���A�<~           �w@                        �-�?&���w�<�            @b@                         �ڦ?����2�<{            �^@������������������������       ��{���<O            �S@������������������������       ����R@1 =,             F@                          s��?�бf[z�<             7@������������������������       �������<             6@������������������������       �      й             �?                          �P�?����X��<�            �m@                        �m��?�;�@�=
             $@������������������������       ���VV���<             @������������������������       ���ܡ�=             @                        �-�?���}j�<�            @l@������������������������       �G8��h��<w            �]@������������������������       ���B��<k            �Z@                         �t�?)��ޔ=             4@                        �[�?�`���<             @                        ��j? ���:&�<             @������������������������       � �A�p�<             @������������������������       �      �             �?������������������������       �      �9             �?        '                  Ʒ�?&���J��<             .@!       $                  9�?�U���]�<              @"       #                 P���?��E.
]�<             @������������������������       ��pV�<              @������������������������       �                     �?%       &                 p۶�?����K�<             @������������������������       �                     �?������������������������       � 0�����<             @(       )                 ��ܵ?5 (�'��<             @������������������������       �                     �?*       +                  `���?
)`����<             @������������������������       �                     �?������������������������       �P�		o<             @-       4                 ��Ѐ?�=��dj�<:             M@.       3                 ���?S�2Ҕ�<	             "@/       0                  �x?�2Y��T�<              @������������������������       ����<             @1       2                 �Yz?��	��>�<             @������������������������       � �e<              @������������������������       �      ҹ             �?������������������������       �      й             �?5       <                 �K��?7�;��]�<1            �H@6       7                  �_�?@]@}u��<             *@������������������������       �D�yT�<             @8       9                  �?��ې���<	             "@������������������������       �p��BjY�<             @:       ;                 0�C�?�*�!��<             @������������������������       �PI=f��<             @������������������������       ��	����<             @=       D                 @8��?�:*�!��<$             B@>       A                 `���?ۼ�"�s�<              @@?       @                 �i�?���?���<             *@������������������������       �t�%*���<             &@������������������������       �  	�;              @B       C                  �/�?Vq8�F�<             3@������������������������       �                     �?������������������������       ��r%1]7�<             2@E       H                 ���?����5�<             @F       G                ��!�?����V�<              @������������������������       �                     �?������������������������       �      �9             �?������������������������       �Xt�'{<              @�t�bh�hhK ��h��R�(KKIKK��h �BH  i���>�4>���'>D�A���>���M�b�9׶���R����A�B#�Vץ	�fٿ *�`UU�?��sUU����UU忭B%X��>)!ʮ�iA>���![P>g8���?XT�d�H�?
�ʱ�`������ֿ�;}�UU�!$�y�#�+��"�l��hWE�ȿA8ݠUU忁�X�E�޽=�������:ʶ�1�?r/
(?�h>��r�[�>  �@��>�~��UU�?*�UU�?���XUU�?&u^LH>�Gգ�a>3���sX��M�$ȍ¿>�kUU�   x�q>�މaUU�?SspUU�?;��͊3L� M_�UU�g|S�*#E>Z�asUU�?BXUU�@����N���3��#h�o܅Z�a�Y��sп5����t��]wUU��N�eUU���,�UU�p�V�Z�B�f`��[���A��?`1��d�N/�[UU�gR� Pm�<K5dUU忣huUU���4"]�%�]����* >�<��?E�T���㿍�A[UU�?>�ڣXE>��[kUU�?�����?(Geod����p�Lt�Ț�wUU�liUU忉�UUU忔t�bubh,h-ubhj)��}�(h9h:hmhnh@Kh;Kh<Kh=G        h?NhGNhDhthAG        h�NhBG        hKh�Kh\Kh�h�KhhK ��h��R�(KK��h��C       �t�bK��R�}�(h@Kh�K+h�hhK ��h��R�(KK+��h��Bh	         &                 �)�?Ɇ�����<�           �}@                        �6Sz?t��ʡ��<�           �|@                        �Ly?�i�&X�<v           `w@                        pF9�??M'��^�<t           @w@                        ���?_z��?X�<q           w@                        pr��?�����<d           @v@������������������������       ��<��n��<[           �u@������������������������       �1]�#���<	             "@	       
                 ��6�?��(�[�<             *@������������������������       �@ ~��<              @������������������������       ���3K?u�<             &@                        �CL?�E�tI�<             @������������������������       �                     �?                        �-�?(������<              @������������������������       �                     �?������������������������       �      ��             �?                        p')�?4�^���<              @������������������������       �                     �?������������������������       �      ��             �?                        `Q�?��N����<U            @U@                         ���?����<6             K@                        `�ռ?��ߐ�b�<             9@                           �?�/T����<             @������������������������       ��5%?	�<             @������������������������       �P���{�<             @������������������������       ���R ��<             3@                         �E�?˟Lo�:�<             =@                        ��\�?�_��r��<             @������������������������       ��H���<�<              @������������������������       �                     �?������������������������       ����ә�<             :@        %                 ��,�?������<             ?@!       $                  ���?��vP�p�<             @"       #                 ��v�?��	GZ�<             @������������������������       �                     �?������������������������       � ��`Up<             @������������������������       �      �             �?������������������������       �	� e��<             8@'       *                 4 �?r(��m��<             *@(       )                 ����?�ܟ��԰<              @������������������������       �                     �?������������������������       �                     �?������������������������       ��U�dތ<             &@�t�bh�hhK ��h��R�(KK+KK��h �BX  ��?` �>�i��"�ƽ��������o3%��w>Z�"�Հ7���,
�4	+��M�iUU�?��~X[W>&�/�UU�?�
��/б?M���c�r��r��UU��g"I,�\��¹dUU忺Z@YUU�r@��8w� -�UU忶Ej\UU��: ��>>��3O>R�Z�X>UU�S";k>F�r_UU�?��eqUU�?%�^UU�?�J��=>�bR@��U�БZUU�?���oUU���V\UU�?��,|�87��`EO��e�|R#��M�n�PzUU�5�XUU�?��UU忱"��@�??n�h��V>  ��X}>��UU�?��vUU�?�2�5��?�t�bubh,h-ubet�b�n_estimators_�K(�init_��sklearn.dummy��DummyClassifier���)��}�(�strategy��prior�hDN�constant�N�	_strategy�jw  �sparse_output_��h�KhLhhK ��h��R�(KK��h��C                      �t�bhTK�class_prior_�hhK ��h��R�(KK��h �C_[4��?	N�<�?��V'�?�t�bh,h-ub�train_score_�hhK ��h��R�(KK(��h �B@  $N���:�?ã�����?�'>�;�?��~��X�?8����Ԡ?4�W �D�?p�P�g�?�F��Yi�?6��=�u?9��Q�bl?�fw>�d?mˡ`r_?�R{�\�R?��ǦM?�h�޿C?�z3��8?���wt1?�_���J)?�����#?_
j��?�L|]?h vg�:?������>��V�%��>а�b\g�>��t7=u�>#hyra�>�Ԓ����>+�XR���>�"�$��>N��G~�>'uC��E�>��)^�>��4=�>�pRP	p�>#h�Q�>��ȵk�{>+�Ưubt>��1�O0k>_�
�c>�t�b�_rng�hth,h-ub��e�memory�NhF�ub.